
module memory_WIDTH8_SIZE8_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13,
         N14, N15, N16, N17, N18, N19, N20, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[7]  ( .D(N13), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N14), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N15), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N16), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N17), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N18), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N19), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N20), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][7]  ( .D(n149), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n148), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n147), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n146), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n145), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n144), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n143), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n142), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n141), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n140), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n139), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n138), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n137), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n136), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n135), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n134), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n133), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n132), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n131), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n130), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n129), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n128), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n127), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n126), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n125), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n124), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n123), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n122), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n121), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n120), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n119), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n118), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n117), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n116), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n115), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n114), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n113), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n112), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n111), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n110), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n109), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n108), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n107), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n106), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n105), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n104), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n103), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n102), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n101), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n100), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n99), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n98), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n97), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n96), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n95), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n94), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n93), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n92), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n91), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n90), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n89), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n88), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n87), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n86), .CK(clk), .Q(\mem[0][0] ) );
  NOR2_X1 U3 ( .A1(n198), .A2(N12), .ZN(n21) );
  BUF_X1 U4 ( .A(N10), .Z(n187) );
  NAND3_X1 U5 ( .A1(N10), .A2(n21), .A3(N11), .ZN(n40) );
  NAND3_X1 U6 ( .A1(N10), .A2(n189), .A3(n58), .ZN(n59) );
  NAND3_X1 U7 ( .A1(N11), .A2(n188), .A3(n58), .ZN(n68) );
  NAND3_X1 U8 ( .A1(N11), .A2(N10), .A3(n58), .ZN(n77) );
  NAND3_X1 U9 ( .A1(n21), .A2(n189), .A3(N10), .ZN(n22) );
  NAND3_X1 U10 ( .A1(n21), .A2(n188), .A3(N11), .ZN(n31) );
  NAND3_X1 U11 ( .A1(n188), .A2(n189), .A3(n58), .ZN(n49) );
  NAND3_X1 U12 ( .A1(n188), .A2(n189), .A3(n21), .ZN(n12) );
  INV_X1 U13 ( .A(wr_en), .ZN(n198) );
  INV_X1 U14 ( .A(N11), .ZN(n189) );
  AND2_X1 U15 ( .A1(N12), .A2(wr_en), .ZN(n58) );
  INV_X1 U16 ( .A(N10), .ZN(n188) );
  OAI21_X1 U17 ( .B1(n12), .B2(n190), .A(n13), .ZN(n86) );
  NAND2_X1 U18 ( .A1(\mem[0][0] ), .A2(n12), .ZN(n13) );
  OAI21_X1 U19 ( .B1(n12), .B2(n191), .A(n14), .ZN(n87) );
  NAND2_X1 U20 ( .A1(\mem[0][1] ), .A2(n12), .ZN(n14) );
  OAI21_X1 U21 ( .B1(n12), .B2(n192), .A(n15), .ZN(n88) );
  NAND2_X1 U22 ( .A1(\mem[0][2] ), .A2(n12), .ZN(n15) );
  OAI21_X1 U23 ( .B1(n12), .B2(n193), .A(n16), .ZN(n89) );
  NAND2_X1 U24 ( .A1(\mem[0][3] ), .A2(n12), .ZN(n16) );
  OAI21_X1 U25 ( .B1(n12), .B2(n194), .A(n17), .ZN(n90) );
  NAND2_X1 U26 ( .A1(\mem[0][4] ), .A2(n12), .ZN(n17) );
  OAI21_X1 U27 ( .B1(n12), .B2(n195), .A(n18), .ZN(n91) );
  NAND2_X1 U28 ( .A1(\mem[0][5] ), .A2(n12), .ZN(n18) );
  OAI21_X1 U29 ( .B1(n12), .B2(n196), .A(n19), .ZN(n92) );
  NAND2_X1 U30 ( .A1(\mem[0][6] ), .A2(n12), .ZN(n19) );
  OAI21_X1 U31 ( .B1(n12), .B2(n197), .A(n20), .ZN(n93) );
  NAND2_X1 U32 ( .A1(\mem[0][7] ), .A2(n12), .ZN(n20) );
  OAI21_X1 U33 ( .B1(n190), .B2(n40), .A(n41), .ZN(n110) );
  NAND2_X1 U34 ( .A1(\mem[3][0] ), .A2(n40), .ZN(n41) );
  OAI21_X1 U35 ( .B1(n191), .B2(n40), .A(n42), .ZN(n111) );
  NAND2_X1 U36 ( .A1(\mem[3][1] ), .A2(n40), .ZN(n42) );
  OAI21_X1 U37 ( .B1(n192), .B2(n40), .A(n43), .ZN(n112) );
  NAND2_X1 U38 ( .A1(\mem[3][2] ), .A2(n40), .ZN(n43) );
  OAI21_X1 U39 ( .B1(n193), .B2(n40), .A(n44), .ZN(n113) );
  NAND2_X1 U40 ( .A1(\mem[3][3] ), .A2(n40), .ZN(n44) );
  OAI21_X1 U41 ( .B1(n194), .B2(n40), .A(n45), .ZN(n114) );
  NAND2_X1 U42 ( .A1(\mem[3][4] ), .A2(n40), .ZN(n45) );
  OAI21_X1 U43 ( .B1(n195), .B2(n40), .A(n46), .ZN(n115) );
  NAND2_X1 U44 ( .A1(\mem[3][5] ), .A2(n40), .ZN(n46) );
  OAI21_X1 U45 ( .B1(n196), .B2(n40), .A(n47), .ZN(n116) );
  NAND2_X1 U46 ( .A1(\mem[3][6] ), .A2(n40), .ZN(n47) );
  OAI21_X1 U47 ( .B1(n197), .B2(n40), .A(n48), .ZN(n117) );
  NAND2_X1 U48 ( .A1(\mem[3][7] ), .A2(n40), .ZN(n48) );
  OAI21_X1 U49 ( .B1(n190), .B2(n59), .A(n60), .ZN(n126) );
  NAND2_X1 U50 ( .A1(\mem[5][0] ), .A2(n59), .ZN(n60) );
  OAI21_X1 U51 ( .B1(n191), .B2(n59), .A(n61), .ZN(n127) );
  NAND2_X1 U52 ( .A1(\mem[5][1] ), .A2(n59), .ZN(n61) );
  OAI21_X1 U53 ( .B1(n192), .B2(n59), .A(n62), .ZN(n128) );
  NAND2_X1 U54 ( .A1(\mem[5][2] ), .A2(n59), .ZN(n62) );
  OAI21_X1 U55 ( .B1(n193), .B2(n59), .A(n63), .ZN(n129) );
  NAND2_X1 U56 ( .A1(\mem[5][3] ), .A2(n59), .ZN(n63) );
  OAI21_X1 U57 ( .B1(n194), .B2(n59), .A(n64), .ZN(n130) );
  NAND2_X1 U58 ( .A1(\mem[5][4] ), .A2(n59), .ZN(n64) );
  OAI21_X1 U59 ( .B1(n195), .B2(n59), .A(n65), .ZN(n131) );
  NAND2_X1 U60 ( .A1(\mem[5][5] ), .A2(n59), .ZN(n65) );
  OAI21_X1 U61 ( .B1(n196), .B2(n59), .A(n66), .ZN(n132) );
  NAND2_X1 U62 ( .A1(\mem[5][6] ), .A2(n59), .ZN(n66) );
  OAI21_X1 U63 ( .B1(n197), .B2(n59), .A(n67), .ZN(n133) );
  NAND2_X1 U64 ( .A1(\mem[5][7] ), .A2(n59), .ZN(n67) );
  OAI21_X1 U65 ( .B1(n190), .B2(n68), .A(n69), .ZN(n134) );
  NAND2_X1 U66 ( .A1(\mem[6][0] ), .A2(n68), .ZN(n69) );
  OAI21_X1 U67 ( .B1(n191), .B2(n68), .A(n70), .ZN(n135) );
  NAND2_X1 U68 ( .A1(\mem[6][1] ), .A2(n68), .ZN(n70) );
  OAI21_X1 U69 ( .B1(n192), .B2(n68), .A(n71), .ZN(n136) );
  NAND2_X1 U70 ( .A1(\mem[6][2] ), .A2(n68), .ZN(n71) );
  OAI21_X1 U71 ( .B1(n193), .B2(n68), .A(n72), .ZN(n137) );
  NAND2_X1 U72 ( .A1(\mem[6][3] ), .A2(n68), .ZN(n72) );
  OAI21_X1 U73 ( .B1(n194), .B2(n68), .A(n73), .ZN(n138) );
  NAND2_X1 U74 ( .A1(\mem[6][4] ), .A2(n68), .ZN(n73) );
  OAI21_X1 U75 ( .B1(n195), .B2(n68), .A(n74), .ZN(n139) );
  NAND2_X1 U76 ( .A1(\mem[6][5] ), .A2(n68), .ZN(n74) );
  OAI21_X1 U77 ( .B1(n196), .B2(n68), .A(n75), .ZN(n140) );
  NAND2_X1 U78 ( .A1(\mem[6][6] ), .A2(n68), .ZN(n75) );
  OAI21_X1 U79 ( .B1(n197), .B2(n68), .A(n76), .ZN(n141) );
  NAND2_X1 U80 ( .A1(\mem[6][7] ), .A2(n68), .ZN(n76) );
  OAI21_X1 U81 ( .B1(n190), .B2(n77), .A(n78), .ZN(n142) );
  NAND2_X1 U82 ( .A1(\mem[7][0] ), .A2(n77), .ZN(n78) );
  OAI21_X1 U83 ( .B1(n191), .B2(n77), .A(n79), .ZN(n143) );
  NAND2_X1 U84 ( .A1(\mem[7][1] ), .A2(n77), .ZN(n79) );
  OAI21_X1 U85 ( .B1(n192), .B2(n77), .A(n80), .ZN(n144) );
  NAND2_X1 U86 ( .A1(\mem[7][2] ), .A2(n77), .ZN(n80) );
  OAI21_X1 U87 ( .B1(n193), .B2(n77), .A(n81), .ZN(n145) );
  NAND2_X1 U88 ( .A1(\mem[7][3] ), .A2(n77), .ZN(n81) );
  OAI21_X1 U89 ( .B1(n194), .B2(n77), .A(n82), .ZN(n146) );
  NAND2_X1 U90 ( .A1(\mem[7][4] ), .A2(n77), .ZN(n82) );
  OAI21_X1 U91 ( .B1(n195), .B2(n77), .A(n83), .ZN(n147) );
  NAND2_X1 U92 ( .A1(\mem[7][5] ), .A2(n77), .ZN(n83) );
  OAI21_X1 U93 ( .B1(n196), .B2(n77), .A(n84), .ZN(n148) );
  NAND2_X1 U94 ( .A1(\mem[7][6] ), .A2(n77), .ZN(n84) );
  OAI21_X1 U95 ( .B1(n197), .B2(n77), .A(n85), .ZN(n149) );
  NAND2_X1 U96 ( .A1(\mem[7][7] ), .A2(n77), .ZN(n85) );
  OAI21_X1 U97 ( .B1(n190), .B2(n22), .A(n23), .ZN(n94) );
  NAND2_X1 U98 ( .A1(\mem[1][0] ), .A2(n22), .ZN(n23) );
  OAI21_X1 U99 ( .B1(n191), .B2(n22), .A(n24), .ZN(n95) );
  NAND2_X1 U100 ( .A1(\mem[1][1] ), .A2(n22), .ZN(n24) );
  OAI21_X1 U101 ( .B1(n192), .B2(n22), .A(n25), .ZN(n96) );
  NAND2_X1 U102 ( .A1(\mem[1][2] ), .A2(n22), .ZN(n25) );
  OAI21_X1 U103 ( .B1(n193), .B2(n22), .A(n26), .ZN(n97) );
  NAND2_X1 U104 ( .A1(\mem[1][3] ), .A2(n22), .ZN(n26) );
  OAI21_X1 U105 ( .B1(n194), .B2(n22), .A(n27), .ZN(n98) );
  NAND2_X1 U106 ( .A1(\mem[1][4] ), .A2(n22), .ZN(n27) );
  OAI21_X1 U107 ( .B1(n195), .B2(n22), .A(n28), .ZN(n99) );
  NAND2_X1 U108 ( .A1(\mem[1][5] ), .A2(n22), .ZN(n28) );
  OAI21_X1 U109 ( .B1(n196), .B2(n22), .A(n29), .ZN(n100) );
  NAND2_X1 U110 ( .A1(\mem[1][6] ), .A2(n22), .ZN(n29) );
  OAI21_X1 U111 ( .B1(n197), .B2(n22), .A(n30), .ZN(n101) );
  NAND2_X1 U112 ( .A1(\mem[1][7] ), .A2(n22), .ZN(n30) );
  OAI21_X1 U113 ( .B1(n190), .B2(n31), .A(n32), .ZN(n102) );
  NAND2_X1 U114 ( .A1(\mem[2][0] ), .A2(n31), .ZN(n32) );
  OAI21_X1 U115 ( .B1(n191), .B2(n31), .A(n33), .ZN(n103) );
  NAND2_X1 U116 ( .A1(\mem[2][1] ), .A2(n31), .ZN(n33) );
  OAI21_X1 U117 ( .B1(n192), .B2(n31), .A(n34), .ZN(n104) );
  NAND2_X1 U118 ( .A1(\mem[2][2] ), .A2(n31), .ZN(n34) );
  OAI21_X1 U119 ( .B1(n193), .B2(n31), .A(n35), .ZN(n105) );
  NAND2_X1 U120 ( .A1(\mem[2][3] ), .A2(n31), .ZN(n35) );
  OAI21_X1 U121 ( .B1(n194), .B2(n31), .A(n36), .ZN(n106) );
  NAND2_X1 U122 ( .A1(\mem[2][4] ), .A2(n31), .ZN(n36) );
  OAI21_X1 U123 ( .B1(n195), .B2(n31), .A(n37), .ZN(n107) );
  NAND2_X1 U124 ( .A1(\mem[2][5] ), .A2(n31), .ZN(n37) );
  OAI21_X1 U125 ( .B1(n196), .B2(n31), .A(n38), .ZN(n108) );
  NAND2_X1 U126 ( .A1(\mem[2][6] ), .A2(n31), .ZN(n38) );
  OAI21_X1 U127 ( .B1(n197), .B2(n31), .A(n39), .ZN(n109) );
  NAND2_X1 U128 ( .A1(\mem[2][7] ), .A2(n31), .ZN(n39) );
  OAI21_X1 U129 ( .B1(n190), .B2(n49), .A(n50), .ZN(n118) );
  NAND2_X1 U130 ( .A1(\mem[4][0] ), .A2(n49), .ZN(n50) );
  OAI21_X1 U131 ( .B1(n191), .B2(n49), .A(n51), .ZN(n119) );
  NAND2_X1 U132 ( .A1(\mem[4][1] ), .A2(n49), .ZN(n51) );
  OAI21_X1 U133 ( .B1(n192), .B2(n49), .A(n52), .ZN(n120) );
  NAND2_X1 U134 ( .A1(\mem[4][2] ), .A2(n49), .ZN(n52) );
  OAI21_X1 U135 ( .B1(n193), .B2(n49), .A(n53), .ZN(n121) );
  NAND2_X1 U136 ( .A1(\mem[4][3] ), .A2(n49), .ZN(n53) );
  OAI21_X1 U137 ( .B1(n194), .B2(n49), .A(n54), .ZN(n122) );
  NAND2_X1 U138 ( .A1(\mem[4][4] ), .A2(n49), .ZN(n54) );
  OAI21_X1 U139 ( .B1(n195), .B2(n49), .A(n55), .ZN(n123) );
  NAND2_X1 U140 ( .A1(\mem[4][5] ), .A2(n49), .ZN(n55) );
  OAI21_X1 U141 ( .B1(n196), .B2(n49), .A(n56), .ZN(n124) );
  NAND2_X1 U142 ( .A1(\mem[4][6] ), .A2(n49), .ZN(n56) );
  OAI21_X1 U143 ( .B1(n197), .B2(n49), .A(n57), .ZN(n125) );
  NAND2_X1 U144 ( .A1(\mem[4][7] ), .A2(n49), .ZN(n57) );
  MUX2_X1 U145 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n1) );
  MUX2_X1 U146 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n2) );
  MUX2_X1 U147 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U148 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U149 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U150 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U151 ( .A(n6), .B(n3), .S(N12), .Z(N20) );
  MUX2_X1 U152 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n7) );
  MUX2_X1 U153 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n8) );
  MUX2_X1 U154 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U155 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n10) );
  MUX2_X1 U156 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n11) );
  MUX2_X1 U157 ( .A(n11), .B(n10), .S(N11), .Z(n150) );
  MUX2_X1 U158 ( .A(n150), .B(n9), .S(N12), .Z(N19) );
  MUX2_X1 U159 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n187), .Z(n151) );
  MUX2_X1 U160 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n187), .Z(n152) );
  MUX2_X1 U161 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U162 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n187), .Z(n154) );
  MUX2_X1 U163 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n187), .Z(n155) );
  MUX2_X1 U164 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U165 ( .A(n156), .B(n153), .S(N12), .Z(N18) );
  MUX2_X1 U166 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n187), .Z(n157) );
  MUX2_X1 U167 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n187), .Z(n158) );
  MUX2_X1 U168 ( .A(n158), .B(n157), .S(N11), .Z(n159) );
  MUX2_X1 U169 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n187), .Z(n160) );
  MUX2_X1 U170 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n187), .Z(n161) );
  MUX2_X1 U171 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U172 ( .A(n162), .B(n159), .S(N12), .Z(N17) );
  MUX2_X1 U173 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n187), .Z(n163) );
  MUX2_X1 U174 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n187), .Z(n164) );
  MUX2_X1 U175 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U176 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n187), .Z(n166) );
  MUX2_X1 U177 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n187), .Z(n167) );
  MUX2_X1 U178 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U179 ( .A(n168), .B(n165), .S(N12), .Z(N16) );
  MUX2_X1 U180 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n169) );
  MUX2_X1 U181 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n187), .Z(n170) );
  MUX2_X1 U182 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U183 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n172) );
  MUX2_X1 U184 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n187), .Z(n173) );
  MUX2_X1 U185 ( .A(n173), .B(n172), .S(N11), .Z(n174) );
  MUX2_X1 U186 ( .A(n174), .B(n171), .S(N12), .Z(N15) );
  MUX2_X1 U187 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n175) );
  MUX2_X1 U188 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n187), .Z(n176) );
  MUX2_X1 U189 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U190 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n178) );
  MUX2_X1 U191 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n187), .Z(n179) );
  MUX2_X1 U192 ( .A(n179), .B(n178), .S(N11), .Z(n180) );
  MUX2_X1 U193 ( .A(n180), .B(n177), .S(N12), .Z(N14) );
  MUX2_X1 U194 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n181) );
  MUX2_X1 U195 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n187), .Z(n182) );
  MUX2_X1 U196 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U197 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n184) );
  MUX2_X1 U198 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n187), .Z(n185) );
  MUX2_X1 U199 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U200 ( .A(n186), .B(n183), .S(N12), .Z(N13) );
  INV_X1 U201 ( .A(data_in[0]), .ZN(n190) );
  INV_X1 U202 ( .A(data_in[1]), .ZN(n191) );
  INV_X1 U203 ( .A(data_in[2]), .ZN(n192) );
  INV_X1 U204 ( .A(data_in[3]), .ZN(n193) );
  INV_X1 U205 ( .A(data_in[4]), .ZN(n194) );
  INV_X1 U206 ( .A(data_in[5]), .ZN(n195) );
  INV_X1 U207 ( .A(data_in[6]), .ZN(n196) );
  INV_X1 U208 ( .A(data_in[7]), .ZN(n197) );
endmodule


module memory_WIDTH8_SIZE64_LOGSIZE6 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [5:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, N15, \mem[63][7] , \mem[63][6] ,
         \mem[63][5] , \mem[63][4] , \mem[63][3] , \mem[63][2] , \mem[63][1] ,
         \mem[63][0] , \mem[62][7] , \mem[62][6] , \mem[62][5] , \mem[62][4] ,
         \mem[62][3] , \mem[62][2] , \mem[62][1] , \mem[62][0] , \mem[61][7] ,
         \mem[61][6] , \mem[61][5] , \mem[61][4] , \mem[61][3] , \mem[61][2] ,
         \mem[61][1] , \mem[61][0] , \mem[60][7] , \mem[60][6] , \mem[60][5] ,
         \mem[60][4] , \mem[60][3] , \mem[60][2] , \mem[60][1] , \mem[60][0] ,
         \mem[59][7] , \mem[59][6] , \mem[59][5] , \mem[59][4] , \mem[59][3] ,
         \mem[59][2] , \mem[59][1] , \mem[59][0] , \mem[58][7] , \mem[58][6] ,
         \mem[58][5] , \mem[58][4] , \mem[58][3] , \mem[58][2] , \mem[58][1] ,
         \mem[58][0] , \mem[57][7] , \mem[57][6] , \mem[57][5] , \mem[57][4] ,
         \mem[57][3] , \mem[57][2] , \mem[57][1] , \mem[57][0] , \mem[56][7] ,
         \mem[56][6] , \mem[56][5] , \mem[56][4] , \mem[56][3] , \mem[56][2] ,
         \mem[56][1] , \mem[56][0] , \mem[55][7] , \mem[55][6] , \mem[55][5] ,
         \mem[55][4] , \mem[55][3] , \mem[55][2] , \mem[55][1] , \mem[55][0] ,
         \mem[54][7] , \mem[54][6] , \mem[54][5] , \mem[54][4] , \mem[54][3] ,
         \mem[54][2] , \mem[54][1] , \mem[54][0] , \mem[53][7] , \mem[53][6] ,
         \mem[53][5] , \mem[53][4] , \mem[53][3] , \mem[53][2] , \mem[53][1] ,
         \mem[53][0] , \mem[52][7] , \mem[52][6] , \mem[52][5] , \mem[52][4] ,
         \mem[52][3] , \mem[52][2] , \mem[52][1] , \mem[52][0] , \mem[51][7] ,
         \mem[51][6] , \mem[51][5] , \mem[51][4] , \mem[51][3] , \mem[51][2] ,
         \mem[51][1] , \mem[51][0] , \mem[50][7] , \mem[50][6] , \mem[50][5] ,
         \mem[50][4] , \mem[50][3] , \mem[50][2] , \mem[50][1] , \mem[50][0] ,
         \mem[49][7] , \mem[49][6] , \mem[49][5] , \mem[49][4] , \mem[49][3] ,
         \mem[49][2] , \mem[49][1] , \mem[49][0] , \mem[48][7] , \mem[48][6] ,
         \mem[48][5] , \mem[48][4] , \mem[48][3] , \mem[48][2] , \mem[48][1] ,
         \mem[48][0] , \mem[47][7] , \mem[47][6] , \mem[47][5] , \mem[47][4] ,
         \mem[47][3] , \mem[47][2] , \mem[47][1] , \mem[47][0] , \mem[46][7] ,
         \mem[46][6] , \mem[46][5] , \mem[46][4] , \mem[46][3] , \mem[46][2] ,
         \mem[46][1] , \mem[46][0] , \mem[45][7] , \mem[45][6] , \mem[45][5] ,
         \mem[45][4] , \mem[45][3] , \mem[45][2] , \mem[45][1] , \mem[45][0] ,
         \mem[44][7] , \mem[44][6] , \mem[44][5] , \mem[44][4] , \mem[44][3] ,
         \mem[44][2] , \mem[44][1] , \mem[44][0] , \mem[43][7] , \mem[43][6] ,
         \mem[43][5] , \mem[43][4] , \mem[43][3] , \mem[43][2] , \mem[43][1] ,
         \mem[43][0] , \mem[42][7] , \mem[42][6] , \mem[42][5] , \mem[42][4] ,
         \mem[42][3] , \mem[42][2] , \mem[42][1] , \mem[42][0] , \mem[41][7] ,
         \mem[41][6] , \mem[41][5] , \mem[41][4] , \mem[41][3] , \mem[41][2] ,
         \mem[41][1] , \mem[41][0] , \mem[40][7] , \mem[40][6] , \mem[40][5] ,
         \mem[40][4] , \mem[40][3] , \mem[40][2] , \mem[40][1] , \mem[40][0] ,
         \mem[39][7] , \mem[39][6] , \mem[39][5] , \mem[39][4] , \mem[39][3] ,
         \mem[39][2] , \mem[39][1] , \mem[39][0] , \mem[38][7] , \mem[38][6] ,
         \mem[38][5] , \mem[38][4] , \mem[38][3] , \mem[38][2] , \mem[38][1] ,
         \mem[38][0] , \mem[37][7] , \mem[37][6] , \mem[37][5] , \mem[37][4] ,
         \mem[37][3] , \mem[37][2] , \mem[37][1] , \mem[37][0] , \mem[36][7] ,
         \mem[36][6] , \mem[36][5] , \mem[36][4] , \mem[36][3] , \mem[36][2] ,
         \mem[36][1] , \mem[36][0] , \mem[35][7] , \mem[35][6] , \mem[35][5] ,
         \mem[35][4] , \mem[35][3] , \mem[35][2] , \mem[35][1] , \mem[35][0] ,
         \mem[34][7] , \mem[34][6] , \mem[34][5] , \mem[34][4] , \mem[34][3] ,
         \mem[34][2] , \mem[34][1] , \mem[34][0] , \mem[33][7] , \mem[33][6] ,
         \mem[33][5] , \mem[33][4] , \mem[33][3] , \mem[33][2] , \mem[33][1] ,
         \mem[33][0] , \mem[32][7] , \mem[32][6] , \mem[32][5] , \mem[32][4] ,
         \mem[32][3] , \mem[32][2] , \mem[32][1] , \mem[32][0] , \mem[31][7] ,
         \mem[31][6] , \mem[31][5] , \mem[31][4] , \mem[31][3] , \mem[31][2] ,
         \mem[31][1] , \mem[31][0] , \mem[30][7] , \mem[30][6] , \mem[30][5] ,
         \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] , \mem[30][0] ,
         \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] , \mem[29][3] ,
         \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[28][7] , \mem[28][6] ,
         \mem[28][5] , \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] ,
         \mem[28][0] , \mem[27][7] , \mem[27][6] , \mem[27][5] , \mem[27][4] ,
         \mem[27][3] , \mem[27][2] , \mem[27][1] , \mem[27][0] , \mem[26][7] ,
         \mem[26][6] , \mem[26][5] , \mem[26][4] , \mem[26][3] , \mem[26][2] ,
         \mem[26][1] , \mem[26][0] , \mem[25][7] , \mem[25][6] , \mem[25][5] ,
         \mem[25][4] , \mem[25][3] , \mem[25][2] , \mem[25][1] , \mem[25][0] ,
         \mem[24][7] , \mem[24][6] , \mem[24][5] , \mem[24][4] , \mem[24][3] ,
         \mem[24][2] , \mem[24][1] , \mem[24][0] , \mem[23][7] , \mem[23][6] ,
         \mem[23][5] , \mem[23][4] , \mem[23][3] , \mem[23][2] , \mem[23][1] ,
         \mem[23][0] , \mem[22][7] , \mem[22][6] , \mem[22][5] , \mem[22][4] ,
         \mem[22][3] , \mem[22][2] , \mem[22][1] , \mem[22][0] , \mem[21][7] ,
         \mem[21][6] , \mem[21][5] , \mem[21][4] , \mem[21][3] , \mem[21][2] ,
         \mem[21][1] , \mem[21][0] , \mem[20][7] , \mem[20][6] , \mem[20][5] ,
         \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] , \mem[20][0] ,
         \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] , \mem[19][3] ,
         \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[18][7] , \mem[18][6] ,
         \mem[18][5] , \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] ,
         \mem[18][0] , \mem[17][7] , \mem[17][6] , \mem[17][5] , \mem[17][4] ,
         \mem[17][3] , \mem[17][2] , \mem[17][1] , \mem[17][0] , \mem[16][7] ,
         \mem[16][6] , \mem[16][5] , \mem[16][4] , \mem[16][3] , \mem[16][2] ,
         \mem[16][1] , \mem[16][0] , \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N19,
         N21, N23, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];
  assign N15 = addr[5];

  DFF_X1 \data_out_reg[4]  ( .D(N19), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[0]  ( .D(N23), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[63][7]  ( .D(n522), .CK(clk), .Q(\mem[63][7] ) );
  DFF_X1 \mem_reg[63][6]  ( .D(n523), .CK(clk), .Q(\mem[63][6] ) );
  DFF_X1 \mem_reg[63][5]  ( .D(n524), .CK(clk), .Q(\mem[63][5] ) );
  DFF_X1 \mem_reg[63][4]  ( .D(n525), .CK(clk), .Q(\mem[63][4] ) );
  DFF_X1 \mem_reg[63][3]  ( .D(n526), .CK(clk), .Q(\mem[63][3] ) );
  DFF_X1 \mem_reg[63][2]  ( .D(n527), .CK(clk), .Q(\mem[63][2] ) );
  DFF_X1 \mem_reg[63][1]  ( .D(n528), .CK(clk), .Q(\mem[63][1] ) );
  DFF_X1 \mem_reg[63][0]  ( .D(n529), .CK(clk), .Q(\mem[63][0] ) );
  DFF_X1 \mem_reg[62][7]  ( .D(n530), .CK(clk), .Q(\mem[62][7] ) );
  DFF_X1 \mem_reg[62][6]  ( .D(n531), .CK(clk), .Q(\mem[62][6] ) );
  DFF_X1 \mem_reg[62][5]  ( .D(n532), .CK(clk), .Q(\mem[62][5] ) );
  DFF_X1 \mem_reg[62][4]  ( .D(n533), .CK(clk), .Q(\mem[62][4] ) );
  DFF_X1 \mem_reg[62][3]  ( .D(n534), .CK(clk), .Q(\mem[62][3] ) );
  DFF_X1 \mem_reg[62][2]  ( .D(n535), .CK(clk), .Q(\mem[62][2] ) );
  DFF_X1 \mem_reg[62][1]  ( .D(n536), .CK(clk), .Q(\mem[62][1] ) );
  DFF_X1 \mem_reg[62][0]  ( .D(n537), .CK(clk), .Q(\mem[62][0] ) );
  DFF_X1 \mem_reg[61][7]  ( .D(n538), .CK(clk), .Q(\mem[61][7] ) );
  DFF_X1 \mem_reg[61][6]  ( .D(n539), .CK(clk), .Q(\mem[61][6] ) );
  DFF_X1 \mem_reg[61][5]  ( .D(n540), .CK(clk), .Q(\mem[61][5] ) );
  DFF_X1 \mem_reg[61][4]  ( .D(n541), .CK(clk), .Q(\mem[61][4] ) );
  DFF_X1 \mem_reg[61][3]  ( .D(n542), .CK(clk), .Q(\mem[61][3] ) );
  DFF_X1 \mem_reg[61][2]  ( .D(n543), .CK(clk), .Q(\mem[61][2] ) );
  DFF_X1 \mem_reg[61][1]  ( .D(n544), .CK(clk), .Q(\mem[61][1] ) );
  DFF_X1 \mem_reg[61][0]  ( .D(n545), .CK(clk), .Q(\mem[61][0] ) );
  DFF_X1 \mem_reg[60][7]  ( .D(n546), .CK(clk), .Q(\mem[60][7] ) );
  DFF_X1 \mem_reg[60][6]  ( .D(n547), .CK(clk), .Q(\mem[60][6] ) );
  DFF_X1 \mem_reg[60][5]  ( .D(n548), .CK(clk), .Q(\mem[60][5] ) );
  DFF_X1 \mem_reg[60][4]  ( .D(n549), .CK(clk), .Q(\mem[60][4] ) );
  DFF_X1 \mem_reg[60][3]  ( .D(n550), .CK(clk), .Q(\mem[60][3] ) );
  DFF_X1 \mem_reg[60][2]  ( .D(n551), .CK(clk), .Q(\mem[60][2] ) );
  DFF_X1 \mem_reg[60][1]  ( .D(n552), .CK(clk), .Q(\mem[60][1] ) );
  DFF_X1 \mem_reg[60][0]  ( .D(n553), .CK(clk), .Q(\mem[60][0] ) );
  DFF_X1 \mem_reg[59][7]  ( .D(n554), .CK(clk), .Q(\mem[59][7] ) );
  DFF_X1 \mem_reg[59][6]  ( .D(n555), .CK(clk), .Q(\mem[59][6] ) );
  DFF_X1 \mem_reg[59][5]  ( .D(n556), .CK(clk), .Q(\mem[59][5] ) );
  DFF_X1 \mem_reg[59][4]  ( .D(n557), .CK(clk), .Q(\mem[59][4] ) );
  DFF_X1 \mem_reg[59][3]  ( .D(n558), .CK(clk), .Q(\mem[59][3] ) );
  DFF_X1 \mem_reg[59][2]  ( .D(n559), .CK(clk), .Q(\mem[59][2] ) );
  DFF_X1 \mem_reg[59][1]  ( .D(n560), .CK(clk), .Q(\mem[59][1] ) );
  DFF_X1 \mem_reg[59][0]  ( .D(n561), .CK(clk), .Q(\mem[59][0] ) );
  DFF_X1 \mem_reg[58][7]  ( .D(n562), .CK(clk), .Q(\mem[58][7] ) );
  DFF_X1 \mem_reg[58][6]  ( .D(n563), .CK(clk), .Q(\mem[58][6] ) );
  DFF_X1 \mem_reg[58][5]  ( .D(n564), .CK(clk), .Q(\mem[58][5] ) );
  DFF_X1 \mem_reg[58][4]  ( .D(n565), .CK(clk), .Q(\mem[58][4] ) );
  DFF_X1 \mem_reg[58][3]  ( .D(n566), .CK(clk), .Q(\mem[58][3] ) );
  DFF_X1 \mem_reg[58][2]  ( .D(n567), .CK(clk), .Q(\mem[58][2] ) );
  DFF_X1 \mem_reg[58][1]  ( .D(n568), .CK(clk), .Q(\mem[58][1] ) );
  DFF_X1 \mem_reg[58][0]  ( .D(n569), .CK(clk), .Q(\mem[58][0] ) );
  DFF_X1 \mem_reg[57][7]  ( .D(n570), .CK(clk), .Q(\mem[57][7] ) );
  DFF_X1 \mem_reg[57][6]  ( .D(n571), .CK(clk), .Q(\mem[57][6] ) );
  DFF_X1 \mem_reg[57][5]  ( .D(n572), .CK(clk), .Q(\mem[57][5] ) );
  DFF_X1 \mem_reg[57][4]  ( .D(n573), .CK(clk), .Q(\mem[57][4] ) );
  DFF_X1 \mem_reg[57][3]  ( .D(n574), .CK(clk), .Q(\mem[57][3] ) );
  DFF_X1 \mem_reg[57][2]  ( .D(n575), .CK(clk), .Q(\mem[57][2] ) );
  DFF_X1 \mem_reg[57][1]  ( .D(n576), .CK(clk), .Q(\mem[57][1] ) );
  DFF_X1 \mem_reg[57][0]  ( .D(n577), .CK(clk), .Q(\mem[57][0] ) );
  DFF_X1 \mem_reg[56][7]  ( .D(n578), .CK(clk), .Q(\mem[56][7] ) );
  DFF_X1 \mem_reg[56][6]  ( .D(n579), .CK(clk), .Q(\mem[56][6] ) );
  DFF_X1 \mem_reg[56][5]  ( .D(n580), .CK(clk), .Q(\mem[56][5] ) );
  DFF_X1 \mem_reg[56][4]  ( .D(n581), .CK(clk), .Q(\mem[56][4] ) );
  DFF_X1 \mem_reg[56][3]  ( .D(n1174), .CK(clk), .Q(\mem[56][3] ) );
  DFF_X1 \mem_reg[56][2]  ( .D(n1175), .CK(clk), .Q(\mem[56][2] ) );
  DFF_X1 \mem_reg[56][1]  ( .D(n1176), .CK(clk), .Q(\mem[56][1] ) );
  DFF_X1 \mem_reg[56][0]  ( .D(n1177), .CK(clk), .Q(\mem[56][0] ) );
  DFF_X1 \mem_reg[55][7]  ( .D(n1178), .CK(clk), .Q(\mem[55][7] ) );
  DFF_X1 \mem_reg[55][6]  ( .D(n1179), .CK(clk), .Q(\mem[55][6] ) );
  DFF_X1 \mem_reg[55][5]  ( .D(n1180), .CK(clk), .Q(\mem[55][5] ) );
  DFF_X1 \mem_reg[55][4]  ( .D(n1181), .CK(clk), .Q(\mem[55][4] ) );
  DFF_X1 \mem_reg[55][3]  ( .D(n1182), .CK(clk), .Q(\mem[55][3] ) );
  DFF_X1 \mem_reg[55][2]  ( .D(n1183), .CK(clk), .Q(\mem[55][2] ) );
  DFF_X1 \mem_reg[55][1]  ( .D(n1184), .CK(clk), .Q(\mem[55][1] ) );
  DFF_X1 \mem_reg[55][0]  ( .D(n1185), .CK(clk), .Q(\mem[55][0] ) );
  DFF_X1 \mem_reg[54][7]  ( .D(n1186), .CK(clk), .Q(\mem[54][7] ) );
  DFF_X1 \mem_reg[54][6]  ( .D(n1187), .CK(clk), .Q(\mem[54][6] ) );
  DFF_X1 \mem_reg[54][5]  ( .D(n1188), .CK(clk), .Q(\mem[54][5] ) );
  DFF_X1 \mem_reg[54][4]  ( .D(n1189), .CK(clk), .Q(\mem[54][4] ) );
  DFF_X1 \mem_reg[54][3]  ( .D(n1190), .CK(clk), .Q(\mem[54][3] ) );
  DFF_X1 \mem_reg[54][2]  ( .D(n1191), .CK(clk), .Q(\mem[54][2] ) );
  DFF_X1 \mem_reg[54][1]  ( .D(n1192), .CK(clk), .Q(\mem[54][1] ) );
  DFF_X1 \mem_reg[54][0]  ( .D(n1193), .CK(clk), .Q(\mem[54][0] ) );
  DFF_X1 \mem_reg[53][7]  ( .D(n1194), .CK(clk), .Q(\mem[53][7] ) );
  DFF_X1 \mem_reg[53][6]  ( .D(n1195), .CK(clk), .Q(\mem[53][6] ) );
  DFF_X1 \mem_reg[53][5]  ( .D(n1196), .CK(clk), .Q(\mem[53][5] ) );
  DFF_X1 \mem_reg[53][4]  ( .D(n1197), .CK(clk), .Q(\mem[53][4] ) );
  DFF_X1 \mem_reg[53][3]  ( .D(n1198), .CK(clk), .Q(\mem[53][3] ) );
  DFF_X1 \mem_reg[53][2]  ( .D(n1199), .CK(clk), .Q(\mem[53][2] ) );
  DFF_X1 \mem_reg[53][1]  ( .D(n1200), .CK(clk), .Q(\mem[53][1] ) );
  DFF_X1 \mem_reg[53][0]  ( .D(n1201), .CK(clk), .Q(\mem[53][0] ) );
  DFF_X1 \mem_reg[52][7]  ( .D(n1202), .CK(clk), .Q(\mem[52][7] ) );
  DFF_X1 \mem_reg[52][6]  ( .D(n1203), .CK(clk), .Q(\mem[52][6] ) );
  DFF_X1 \mem_reg[52][5]  ( .D(n1204), .CK(clk), .Q(\mem[52][5] ) );
  DFF_X1 \mem_reg[52][4]  ( .D(n1205), .CK(clk), .Q(\mem[52][4] ) );
  DFF_X1 \mem_reg[52][3]  ( .D(n1206), .CK(clk), .Q(\mem[52][3] ) );
  DFF_X1 \mem_reg[52][2]  ( .D(n1207), .CK(clk), .Q(\mem[52][2] ) );
  DFF_X1 \mem_reg[52][1]  ( .D(n1208), .CK(clk), .Q(\mem[52][1] ) );
  DFF_X1 \mem_reg[52][0]  ( .D(n1209), .CK(clk), .Q(\mem[52][0] ) );
  DFF_X1 \mem_reg[51][7]  ( .D(n1210), .CK(clk), .Q(\mem[51][7] ) );
  DFF_X1 \mem_reg[51][6]  ( .D(n1211), .CK(clk), .Q(\mem[51][6] ) );
  DFF_X1 \mem_reg[51][5]  ( .D(n1212), .CK(clk), .Q(\mem[51][5] ) );
  DFF_X1 \mem_reg[51][4]  ( .D(n1213), .CK(clk), .Q(\mem[51][4] ) );
  DFF_X1 \mem_reg[51][3]  ( .D(n1214), .CK(clk), .Q(\mem[51][3] ) );
  DFF_X1 \mem_reg[51][2]  ( .D(n1215), .CK(clk), .Q(\mem[51][2] ) );
  DFF_X1 \mem_reg[51][1]  ( .D(n1216), .CK(clk), .Q(\mem[51][1] ) );
  DFF_X1 \mem_reg[51][0]  ( .D(n1217), .CK(clk), .Q(\mem[51][0] ) );
  DFF_X1 \mem_reg[50][7]  ( .D(n1218), .CK(clk), .Q(\mem[50][7] ) );
  DFF_X1 \mem_reg[50][6]  ( .D(n1219), .CK(clk), .Q(\mem[50][6] ) );
  DFF_X1 \mem_reg[50][5]  ( .D(n1220), .CK(clk), .Q(\mem[50][5] ) );
  DFF_X1 \mem_reg[50][4]  ( .D(n1221), .CK(clk), .Q(\mem[50][4] ) );
  DFF_X1 \mem_reg[50][3]  ( .D(n1222), .CK(clk), .Q(\mem[50][3] ) );
  DFF_X1 \mem_reg[50][2]  ( .D(n1223), .CK(clk), .Q(\mem[50][2] ) );
  DFF_X1 \mem_reg[50][1]  ( .D(n1224), .CK(clk), .Q(\mem[50][1] ) );
  DFF_X1 \mem_reg[50][0]  ( .D(n1225), .CK(clk), .Q(\mem[50][0] ) );
  DFF_X1 \mem_reg[49][7]  ( .D(n1226), .CK(clk), .Q(\mem[49][7] ) );
  DFF_X1 \mem_reg[49][6]  ( .D(n1227), .CK(clk), .Q(\mem[49][6] ) );
  DFF_X1 \mem_reg[49][5]  ( .D(n1228), .CK(clk), .Q(\mem[49][5] ) );
  DFF_X1 \mem_reg[49][4]  ( .D(n1229), .CK(clk), .Q(\mem[49][4] ) );
  DFF_X1 \mem_reg[49][3]  ( .D(n1230), .CK(clk), .Q(\mem[49][3] ) );
  DFF_X1 \mem_reg[49][2]  ( .D(n1231), .CK(clk), .Q(\mem[49][2] ) );
  DFF_X1 \mem_reg[49][1]  ( .D(n1232), .CK(clk), .Q(\mem[49][1] ) );
  DFF_X1 \mem_reg[49][0]  ( .D(n1233), .CK(clk), .Q(\mem[49][0] ) );
  DFF_X1 \mem_reg[48][7]  ( .D(n1234), .CK(clk), .Q(\mem[48][7] ) );
  DFF_X1 \mem_reg[48][6]  ( .D(n1235), .CK(clk), .Q(\mem[48][6] ) );
  DFF_X1 \mem_reg[48][5]  ( .D(n1236), .CK(clk), .Q(\mem[48][5] ) );
  DFF_X1 \mem_reg[48][4]  ( .D(n1237), .CK(clk), .Q(\mem[48][4] ) );
  DFF_X1 \mem_reg[48][3]  ( .D(n1238), .CK(clk), .Q(\mem[48][3] ) );
  DFF_X1 \mem_reg[48][2]  ( .D(n1239), .CK(clk), .Q(\mem[48][2] ) );
  DFF_X1 \mem_reg[48][1]  ( .D(n1240), .CK(clk), .Q(\mem[48][1] ) );
  DFF_X1 \mem_reg[48][0]  ( .D(n1241), .CK(clk), .Q(\mem[48][0] ) );
  DFF_X1 \mem_reg[47][7]  ( .D(n1242), .CK(clk), .Q(\mem[47][7] ) );
  DFF_X1 \mem_reg[47][6]  ( .D(n1243), .CK(clk), .Q(\mem[47][6] ) );
  DFF_X1 \mem_reg[47][5]  ( .D(n1244), .CK(clk), .Q(\mem[47][5] ) );
  DFF_X1 \mem_reg[47][4]  ( .D(n1245), .CK(clk), .Q(\mem[47][4] ) );
  DFF_X1 \mem_reg[47][3]  ( .D(n1246), .CK(clk), .Q(\mem[47][3] ) );
  DFF_X1 \mem_reg[47][2]  ( .D(n1247), .CK(clk), .Q(\mem[47][2] ) );
  DFF_X1 \mem_reg[47][1]  ( .D(n1248), .CK(clk), .Q(\mem[47][1] ) );
  DFF_X1 \mem_reg[47][0]  ( .D(n1249), .CK(clk), .Q(\mem[47][0] ) );
  DFF_X1 \mem_reg[46][7]  ( .D(n1250), .CK(clk), .Q(\mem[46][7] ) );
  DFF_X1 \mem_reg[46][6]  ( .D(n1251), .CK(clk), .Q(\mem[46][6] ) );
  DFF_X1 \mem_reg[46][5]  ( .D(n1252), .CK(clk), .Q(\mem[46][5] ) );
  DFF_X1 \mem_reg[46][4]  ( .D(n1253), .CK(clk), .Q(\mem[46][4] ) );
  DFF_X1 \mem_reg[46][3]  ( .D(n1254), .CK(clk), .Q(\mem[46][3] ) );
  DFF_X1 \mem_reg[46][2]  ( .D(n1255), .CK(clk), .Q(\mem[46][2] ) );
  DFF_X1 \mem_reg[46][1]  ( .D(n1256), .CK(clk), .Q(\mem[46][1] ) );
  DFF_X1 \mem_reg[46][0]  ( .D(n1257), .CK(clk), .Q(\mem[46][0] ) );
  DFF_X1 \mem_reg[45][7]  ( .D(n1258), .CK(clk), .Q(\mem[45][7] ) );
  DFF_X1 \mem_reg[45][6]  ( .D(n1259), .CK(clk), .Q(\mem[45][6] ) );
  DFF_X1 \mem_reg[45][5]  ( .D(n1260), .CK(clk), .Q(\mem[45][5] ) );
  DFF_X1 \mem_reg[45][4]  ( .D(n1261), .CK(clk), .Q(\mem[45][4] ) );
  DFF_X1 \mem_reg[45][3]  ( .D(n1262), .CK(clk), .Q(\mem[45][3] ) );
  DFF_X1 \mem_reg[45][2]  ( .D(n1263), .CK(clk), .Q(\mem[45][2] ) );
  DFF_X1 \mem_reg[45][1]  ( .D(n1264), .CK(clk), .Q(\mem[45][1] ) );
  DFF_X1 \mem_reg[45][0]  ( .D(n1265), .CK(clk), .Q(\mem[45][0] ) );
  DFF_X1 \mem_reg[44][7]  ( .D(n1266), .CK(clk), .Q(\mem[44][7] ) );
  DFF_X1 \mem_reg[44][6]  ( .D(n1267), .CK(clk), .Q(\mem[44][6] ) );
  DFF_X1 \mem_reg[44][5]  ( .D(n1268), .CK(clk), .Q(\mem[44][5] ) );
  DFF_X1 \mem_reg[44][4]  ( .D(n1269), .CK(clk), .Q(\mem[44][4] ) );
  DFF_X1 \mem_reg[44][3]  ( .D(n1270), .CK(clk), .Q(\mem[44][3] ) );
  DFF_X1 \mem_reg[44][2]  ( .D(n1271), .CK(clk), .Q(\mem[44][2] ) );
  DFF_X1 \mem_reg[44][1]  ( .D(n1272), .CK(clk), .Q(\mem[44][1] ) );
  DFF_X1 \mem_reg[44][0]  ( .D(n1273), .CK(clk), .Q(\mem[44][0] ) );
  DFF_X1 \mem_reg[43][7]  ( .D(n1274), .CK(clk), .Q(\mem[43][7] ) );
  DFF_X1 \mem_reg[43][6]  ( .D(n1275), .CK(clk), .Q(\mem[43][6] ) );
  DFF_X1 \mem_reg[43][5]  ( .D(n1276), .CK(clk), .Q(\mem[43][5] ) );
  DFF_X1 \mem_reg[43][4]  ( .D(n1277), .CK(clk), .Q(\mem[43][4] ) );
  DFF_X1 \mem_reg[43][3]  ( .D(n1278), .CK(clk), .Q(\mem[43][3] ) );
  DFF_X1 \mem_reg[43][2]  ( .D(n1279), .CK(clk), .Q(\mem[43][2] ) );
  DFF_X1 \mem_reg[43][1]  ( .D(n1280), .CK(clk), .Q(\mem[43][1] ) );
  DFF_X1 \mem_reg[43][0]  ( .D(n1281), .CK(clk), .Q(\mem[43][0] ) );
  DFF_X1 \mem_reg[42][7]  ( .D(n1282), .CK(clk), .Q(\mem[42][7] ) );
  DFF_X1 \mem_reg[42][6]  ( .D(n1283), .CK(clk), .Q(\mem[42][6] ) );
  DFF_X1 \mem_reg[42][5]  ( .D(n1284), .CK(clk), .Q(\mem[42][5] ) );
  DFF_X1 \mem_reg[42][4]  ( .D(n1285), .CK(clk), .Q(\mem[42][4] ) );
  DFF_X1 \mem_reg[42][3]  ( .D(n1286), .CK(clk), .Q(\mem[42][3] ) );
  DFF_X1 \mem_reg[42][2]  ( .D(n1287), .CK(clk), .Q(\mem[42][2] ) );
  DFF_X1 \mem_reg[42][1]  ( .D(n1288), .CK(clk), .Q(\mem[42][1] ) );
  DFF_X1 \mem_reg[42][0]  ( .D(n1289), .CK(clk), .Q(\mem[42][0] ) );
  DFF_X1 \mem_reg[41][7]  ( .D(n1290), .CK(clk), .Q(\mem[41][7] ) );
  DFF_X1 \mem_reg[41][6]  ( .D(n1291), .CK(clk), .Q(\mem[41][6] ) );
  DFF_X1 \mem_reg[41][5]  ( .D(n1292), .CK(clk), .Q(\mem[41][5] ) );
  DFF_X1 \mem_reg[41][4]  ( .D(n1293), .CK(clk), .Q(\mem[41][4] ) );
  DFF_X1 \mem_reg[41][3]  ( .D(n1294), .CK(clk), .Q(\mem[41][3] ) );
  DFF_X1 \mem_reg[41][2]  ( .D(n1295), .CK(clk), .Q(\mem[41][2] ) );
  DFF_X1 \mem_reg[41][1]  ( .D(n1296), .CK(clk), .Q(\mem[41][1] ) );
  DFF_X1 \mem_reg[41][0]  ( .D(n1297), .CK(clk), .Q(\mem[41][0] ) );
  DFF_X1 \mem_reg[40][7]  ( .D(n1298), .CK(clk), .Q(\mem[40][7] ) );
  DFF_X1 \mem_reg[40][6]  ( .D(n1299), .CK(clk), .Q(\mem[40][6] ) );
  DFF_X1 \mem_reg[40][5]  ( .D(n1300), .CK(clk), .Q(\mem[40][5] ) );
  DFF_X1 \mem_reg[40][4]  ( .D(n1301), .CK(clk), .Q(\mem[40][4] ) );
  DFF_X1 \mem_reg[40][3]  ( .D(n1302), .CK(clk), .Q(\mem[40][3] ) );
  DFF_X1 \mem_reg[40][2]  ( .D(n1303), .CK(clk), .Q(\mem[40][2] ) );
  DFF_X1 \mem_reg[40][1]  ( .D(n1304), .CK(clk), .Q(\mem[40][1] ) );
  DFF_X1 \mem_reg[40][0]  ( .D(n1305), .CK(clk), .Q(\mem[40][0] ) );
  DFF_X1 \mem_reg[39][7]  ( .D(n1306), .CK(clk), .Q(\mem[39][7] ) );
  DFF_X1 \mem_reg[39][6]  ( .D(n1307), .CK(clk), .Q(\mem[39][6] ) );
  DFF_X1 \mem_reg[39][5]  ( .D(n1308), .CK(clk), .Q(\mem[39][5] ) );
  DFF_X1 \mem_reg[39][4]  ( .D(n1309), .CK(clk), .Q(\mem[39][4] ) );
  DFF_X1 \mem_reg[39][3]  ( .D(n1310), .CK(clk), .Q(\mem[39][3] ) );
  DFF_X1 \mem_reg[39][2]  ( .D(n1311), .CK(clk), .Q(\mem[39][2] ) );
  DFF_X1 \mem_reg[39][1]  ( .D(n1312), .CK(clk), .Q(\mem[39][1] ) );
  DFF_X1 \mem_reg[39][0]  ( .D(n1313), .CK(clk), .Q(\mem[39][0] ) );
  DFF_X1 \mem_reg[38][7]  ( .D(n1314), .CK(clk), .Q(\mem[38][7] ) );
  DFF_X1 \mem_reg[38][6]  ( .D(n1315), .CK(clk), .Q(\mem[38][6] ) );
  DFF_X1 \mem_reg[38][5]  ( .D(n1316), .CK(clk), .Q(\mem[38][5] ) );
  DFF_X1 \mem_reg[38][4]  ( .D(n1317), .CK(clk), .Q(\mem[38][4] ) );
  DFF_X1 \mem_reg[38][3]  ( .D(n1318), .CK(clk), .Q(\mem[38][3] ) );
  DFF_X1 \mem_reg[38][2]  ( .D(n1319), .CK(clk), .Q(\mem[38][2] ) );
  DFF_X1 \mem_reg[38][1]  ( .D(n1320), .CK(clk), .Q(\mem[38][1] ) );
  DFF_X1 \mem_reg[38][0]  ( .D(n1321), .CK(clk), .Q(\mem[38][0] ) );
  DFF_X1 \mem_reg[37][7]  ( .D(n1322), .CK(clk), .Q(\mem[37][7] ) );
  DFF_X1 \mem_reg[37][6]  ( .D(n1323), .CK(clk), .Q(\mem[37][6] ) );
  DFF_X1 \mem_reg[37][5]  ( .D(n1324), .CK(clk), .Q(\mem[37][5] ) );
  DFF_X1 \mem_reg[37][4]  ( .D(n1325), .CK(clk), .Q(\mem[37][4] ) );
  DFF_X1 \mem_reg[37][3]  ( .D(n1326), .CK(clk), .Q(\mem[37][3] ) );
  DFF_X1 \mem_reg[37][2]  ( .D(n1327), .CK(clk), .Q(\mem[37][2] ) );
  DFF_X1 \mem_reg[37][1]  ( .D(n1328), .CK(clk), .Q(\mem[37][1] ) );
  DFF_X1 \mem_reg[37][0]  ( .D(n1329), .CK(clk), .Q(\mem[37][0] ) );
  DFF_X1 \mem_reg[36][7]  ( .D(n1330), .CK(clk), .Q(\mem[36][7] ) );
  DFF_X1 \mem_reg[36][6]  ( .D(n1331), .CK(clk), .Q(\mem[36][6] ) );
  DFF_X1 \mem_reg[36][5]  ( .D(n1332), .CK(clk), .Q(\mem[36][5] ) );
  DFF_X1 \mem_reg[36][4]  ( .D(n1333), .CK(clk), .Q(\mem[36][4] ) );
  DFF_X1 \mem_reg[36][3]  ( .D(n1334), .CK(clk), .Q(\mem[36][3] ) );
  DFF_X1 \mem_reg[36][2]  ( .D(n1335), .CK(clk), .Q(\mem[36][2] ) );
  DFF_X1 \mem_reg[36][1]  ( .D(n1336), .CK(clk), .Q(\mem[36][1] ) );
  DFF_X1 \mem_reg[36][0]  ( .D(n1337), .CK(clk), .Q(\mem[36][0] ) );
  DFF_X1 \mem_reg[35][7]  ( .D(n1338), .CK(clk), .Q(\mem[35][7] ) );
  DFF_X1 \mem_reg[35][6]  ( .D(n1339), .CK(clk), .Q(\mem[35][6] ) );
  DFF_X1 \mem_reg[35][5]  ( .D(n1340), .CK(clk), .Q(\mem[35][5] ) );
  DFF_X1 \mem_reg[35][4]  ( .D(n1341), .CK(clk), .Q(\mem[35][4] ) );
  DFF_X1 \mem_reg[35][3]  ( .D(n1342), .CK(clk), .Q(\mem[35][3] ) );
  DFF_X1 \mem_reg[35][2]  ( .D(n1343), .CK(clk), .Q(\mem[35][2] ) );
  DFF_X1 \mem_reg[35][1]  ( .D(n1344), .CK(clk), .Q(\mem[35][1] ) );
  DFF_X1 \mem_reg[35][0]  ( .D(n1345), .CK(clk), .Q(\mem[35][0] ) );
  DFF_X1 \mem_reg[34][7]  ( .D(n1346), .CK(clk), .Q(\mem[34][7] ) );
  DFF_X1 \mem_reg[34][6]  ( .D(n1347), .CK(clk), .Q(\mem[34][6] ) );
  DFF_X1 \mem_reg[34][5]  ( .D(n1348), .CK(clk), .Q(\mem[34][5] ) );
  DFF_X1 \mem_reg[34][4]  ( .D(n1349), .CK(clk), .Q(\mem[34][4] ) );
  DFF_X1 \mem_reg[34][3]  ( .D(n1350), .CK(clk), .Q(\mem[34][3] ) );
  DFF_X1 \mem_reg[34][2]  ( .D(n1351), .CK(clk), .Q(\mem[34][2] ) );
  DFF_X1 \mem_reg[34][1]  ( .D(n1352), .CK(clk), .Q(\mem[34][1] ) );
  DFF_X1 \mem_reg[34][0]  ( .D(n1353), .CK(clk), .Q(\mem[34][0] ) );
  DFF_X1 \mem_reg[33][7]  ( .D(n1354), .CK(clk), .Q(\mem[33][7] ) );
  DFF_X1 \mem_reg[33][6]  ( .D(n1355), .CK(clk), .Q(\mem[33][6] ) );
  DFF_X1 \mem_reg[33][5]  ( .D(n1356), .CK(clk), .Q(\mem[33][5] ) );
  DFF_X1 \mem_reg[33][4]  ( .D(n1357), .CK(clk), .Q(\mem[33][4] ) );
  DFF_X1 \mem_reg[33][3]  ( .D(n1358), .CK(clk), .Q(\mem[33][3] ) );
  DFF_X1 \mem_reg[33][2]  ( .D(n1359), .CK(clk), .Q(\mem[33][2] ) );
  DFF_X1 \mem_reg[33][1]  ( .D(n1360), .CK(clk), .Q(\mem[33][1] ) );
  DFF_X1 \mem_reg[33][0]  ( .D(n1361), .CK(clk), .Q(\mem[33][0] ) );
  DFF_X1 \mem_reg[32][7]  ( .D(n1362), .CK(clk), .Q(\mem[32][7] ) );
  DFF_X1 \mem_reg[32][6]  ( .D(n1363), .CK(clk), .Q(\mem[32][6] ) );
  DFF_X1 \mem_reg[32][5]  ( .D(n1364), .CK(clk), .Q(\mem[32][5] ) );
  DFF_X1 \mem_reg[32][4]  ( .D(n1365), .CK(clk), .Q(\mem[32][4] ) );
  DFF_X1 \mem_reg[32][3]  ( .D(n1366), .CK(clk), .Q(\mem[32][3] ) );
  DFF_X1 \mem_reg[32][2]  ( .D(n1367), .CK(clk), .Q(\mem[32][2] ) );
  DFF_X1 \mem_reg[32][1]  ( .D(n1368), .CK(clk), .Q(\mem[32][1] ) );
  DFF_X1 \mem_reg[32][0]  ( .D(n1369), .CK(clk), .Q(\mem[32][0] ) );
  DFF_X1 \mem_reg[31][7]  ( .D(n1370), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n1371), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n1372), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n1373), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n1374), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n1375), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n1376), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n1377), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n1378), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n1379), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n1380), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n1381), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n1382), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n1383), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n1384), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n1385), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n1386), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n1387), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n1388), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n1389), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n1390), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n1391), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n1392), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n1393), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n1394), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n1395), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n1396), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n1397), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n1398), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n1399), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n1400), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n1401), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n1402), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n1403), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n1404), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n1405), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n1406), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n1407), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n1408), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n1409), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n1410), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n1411), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n1412), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n1413), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n1414), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n1415), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n1416), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n1417), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n1418), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n1419), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n1420), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n1421), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n1422), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n1423), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n1424), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n1425), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n1426), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n1427), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n1428), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n1429), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n1430), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n1431), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n1432), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n1433), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n1434), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n1435), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n1436), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n1437), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n1438), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n1439), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n1440), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n1441), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n1442), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n1443), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n1444), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n1445), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n1446), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n1447), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n1448), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n1449), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n1450), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n1451), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n1452), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n1453), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n1454), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n1455), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n1456), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n1457), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n1458), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n1459), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n1460), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n1461), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n1462), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n1463), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n1464), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n1465), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n1466), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n1467), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n1468), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n1469), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n1470), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n1471), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n1472), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n1473), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n1474), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n1475), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n1476), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n1477), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n1478), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n1479), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n1480), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n1481), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n1482), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n1483), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n1484), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n1485), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n1486), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n1487), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n1488), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n1489), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n1490), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n1491), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n1492), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n1493), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n1494), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n1495), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n1496), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n1497), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n1498), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n1499), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n1500), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n1501), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n1502), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n1503), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n1504), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n1505), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n1506), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n1507), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n1508), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n1509), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n1510), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n1511), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n1512), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n1513), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n1514), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n1515), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n1516), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n1517), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n1518), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n1519), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n1520), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n1521), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n1522), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n1523), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n1524), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n1525), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n1526), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n1527), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n1528), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n1529), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n1530), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n1531), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n1532), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n1533), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n1534), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n1535), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n1536), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n1537), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n1538), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n1539), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n1540), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n1541), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n1542), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n1543), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n1544), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n1545), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n1546), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n1547), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n1548), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n1549), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n1550), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n1551), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n1552), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n1553), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n1554), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n1555), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n1556), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n1557), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n1558), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n1559), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n1560), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n1561), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n1562), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n1563), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n1564), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n1565), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n1566), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n1567), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n1568), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n1569), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n1570), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n1571), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n1572), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n1573), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n1574), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n1575), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n1576), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n1577), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n1578), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n1579), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n1580), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n1581), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n1582), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n1583), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n1584), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n1585), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n1586), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n1587), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n1588), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n1589), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n1590), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n1591), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n1592), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n1593), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n1594), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n1595), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n1596), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n1597), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n1598), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n1599), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n1600), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n1601), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n1602), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n1603), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n1604), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n1605), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n1606), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n1607), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n1608), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n1609), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n1610), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n1611), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n1612), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n1613), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n1614), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n1615), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n1616), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n1617), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n1618), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n1619), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n1620), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n1621), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n1622), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n1623), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n1624), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n1625), .CK(clk), .Q(\mem[0][0] ) );
  NOR3_X2 U523 ( .A1(N11), .A2(N12), .A3(n510), .ZN(n591) );
  NOR3_X2 U533 ( .A1(N11), .A2(N12), .A3(n518), .ZN(n602) );
  NOR3_X2 U543 ( .A1(n510), .A2(N12), .A3(n519), .ZN(n612) );
  NOR3_X2 U553 ( .A1(n518), .A2(N12), .A3(n519), .ZN(n622) );
  DFF_X1 \data_out_reg[2]  ( .D(N21), .CK(clk), .Q(data_out[2]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n219), .SI(n250), .SE(n1690), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n343), .SI(n374), .SE(n1690), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n95), .SI(n126), .SE(n1690), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n405), .SI(n436), .SE(n1690), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n467), .SI(n498), .SE(n1690), .CK(clk), .Q(
        data_out[7]) );
  BUF_X2 U3 ( .A(N10), .Z(n513) );
  BUF_X1 U4 ( .A(N12), .Z(n501) );
  BUF_X1 U5 ( .A(N11), .Z(n503) );
  CLKBUF_X1 U6 ( .A(N11), .Z(n509) );
  AND3_X1 U7 ( .A1(N10), .A2(n519), .A3(N12), .ZN(n642) );
  AND3_X1 U8 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n662) );
  CLKBUF_X3 U9 ( .A(N10), .Z(n510) );
  CLKBUF_X3 U10 ( .A(N10), .Z(n511) );
  CLKBUF_X2 U11 ( .A(N10), .Z(n512) );
  BUF_X1 U12 ( .A(n516), .Z(n1) );
  AND4_X1 U13 ( .A1(N13), .A2(wr_en), .A3(n521), .A4(n1690), .ZN(n672) );
  AND4_X1 U14 ( .A1(N14), .A2(wr_en), .A3(n520), .A4(n1690), .ZN(n745) );
  AND4_X1 U15 ( .A1(N14), .A2(N13), .A3(wr_en), .A4(n1690), .ZN(n818) );
  AND4_X1 U16 ( .A1(N15), .A2(wr_en), .A3(n520), .A4(n521), .ZN(n891) );
  AND4_X1 U17 ( .A1(N15), .A2(N13), .A3(wr_en), .A4(n521), .ZN(n964) );
  AND4_X1 U18 ( .A1(N15), .A2(N14), .A3(wr_en), .A4(n520), .ZN(n1037) );
  AND4_X1 U19 ( .A1(N15), .A2(N14), .A3(N13), .A4(wr_en), .ZN(n1110) );
  BUF_X1 U20 ( .A(n516), .Z(n515) );
  BUF_X1 U21 ( .A(n516), .Z(n514) );
  BUF_X1 U22 ( .A(N10), .Z(n516) );
  BUF_X1 U23 ( .A(n509), .Z(n507) );
  BUF_X1 U24 ( .A(n509), .Z(n508) );
  BUF_X1 U25 ( .A(n509), .Z(n506) );
  BUF_X1 U26 ( .A(N11), .Z(n504) );
  BUF_X1 U27 ( .A(n509), .Z(n505) );
  INV_X1 U28 ( .A(n594), .ZN(n1688) );
  INV_X1 U29 ( .A(n604), .ZN(n1687) );
  INV_X1 U30 ( .A(n614), .ZN(n1686) );
  INV_X1 U31 ( .A(n664), .ZN(n1681) );
  INV_X1 U32 ( .A(n674), .ZN(n1680) );
  INV_X1 U33 ( .A(n683), .ZN(n1679) );
  INV_X1 U34 ( .A(n692), .ZN(n1678) );
  INV_X1 U35 ( .A(n737), .ZN(n1673) );
  INV_X1 U36 ( .A(n747), .ZN(n1672) );
  INV_X1 U37 ( .A(n756), .ZN(n1671) );
  INV_X1 U38 ( .A(n765), .ZN(n1670) );
  INV_X1 U39 ( .A(n810), .ZN(n1665) );
  INV_X1 U40 ( .A(n820), .ZN(n1664) );
  INV_X1 U41 ( .A(n829), .ZN(n1663) );
  INV_X1 U42 ( .A(n838), .ZN(n1662) );
  INV_X1 U43 ( .A(n883), .ZN(n1657) );
  INV_X1 U44 ( .A(n893), .ZN(n1656) );
  INV_X1 U45 ( .A(n902), .ZN(n1655) );
  INV_X1 U46 ( .A(n911), .ZN(n1654) );
  INV_X1 U47 ( .A(n956), .ZN(n1649) );
  INV_X1 U48 ( .A(n966), .ZN(n1648) );
  INV_X1 U49 ( .A(n975), .ZN(n1647) );
  INV_X1 U50 ( .A(n984), .ZN(n1646) );
  INV_X1 U51 ( .A(n1029), .ZN(n1641) );
  INV_X1 U52 ( .A(n1039), .ZN(n1640) );
  INV_X1 U53 ( .A(n1048), .ZN(n1639) );
  INV_X1 U54 ( .A(n1057), .ZN(n1638) );
  INV_X1 U55 ( .A(n1102), .ZN(n1633) );
  INV_X1 U56 ( .A(n1112), .ZN(n1632) );
  INV_X1 U57 ( .A(n1121), .ZN(n1631) );
  INV_X1 U58 ( .A(n1130), .ZN(n1630) );
  INV_X1 U59 ( .A(n624), .ZN(n1685) );
  INV_X1 U60 ( .A(n634), .ZN(n1684) );
  INV_X1 U61 ( .A(n644), .ZN(n1683) );
  INV_X1 U62 ( .A(n654), .ZN(n1682) );
  INV_X1 U63 ( .A(n701), .ZN(n1677) );
  INV_X1 U64 ( .A(n710), .ZN(n1676) );
  INV_X1 U65 ( .A(n719), .ZN(n1675) );
  INV_X1 U66 ( .A(n728), .ZN(n1674) );
  INV_X1 U67 ( .A(n774), .ZN(n1669) );
  INV_X1 U68 ( .A(n783), .ZN(n1668) );
  INV_X1 U69 ( .A(n792), .ZN(n1667) );
  INV_X1 U70 ( .A(n801), .ZN(n1666) );
  INV_X1 U71 ( .A(n847), .ZN(n1661) );
  INV_X1 U72 ( .A(n856), .ZN(n1660) );
  INV_X1 U73 ( .A(n865), .ZN(n1659) );
  INV_X1 U74 ( .A(n874), .ZN(n1658) );
  INV_X1 U75 ( .A(n920), .ZN(n1653) );
  INV_X1 U76 ( .A(n929), .ZN(n1652) );
  INV_X1 U77 ( .A(n938), .ZN(n1651) );
  INV_X1 U78 ( .A(n947), .ZN(n1650) );
  INV_X1 U79 ( .A(n993), .ZN(n1645) );
  INV_X1 U80 ( .A(n1002), .ZN(n1644) );
  INV_X1 U81 ( .A(n1011), .ZN(n1643) );
  INV_X1 U82 ( .A(n1020), .ZN(n1642) );
  INV_X1 U83 ( .A(n1066), .ZN(n1637) );
  INV_X1 U84 ( .A(n1075), .ZN(n1636) );
  INV_X1 U85 ( .A(n1084), .ZN(n1635) );
  INV_X1 U86 ( .A(n1093), .ZN(n1634) );
  INV_X1 U87 ( .A(n1139), .ZN(n1629) );
  INV_X1 U88 ( .A(n1148), .ZN(n1628) );
  INV_X1 U89 ( .A(n1157), .ZN(n1627) );
  INV_X1 U90 ( .A(n1166), .ZN(n1626) );
  INV_X1 U91 ( .A(n583), .ZN(n1689) );
  BUF_X1 U92 ( .A(N13), .Z(n499) );
  NAND2_X1 U93 ( .A1(n591), .A2(n592), .ZN(n583) );
  NAND2_X1 U94 ( .A1(n602), .A2(n592), .ZN(n594) );
  NAND2_X1 U95 ( .A1(n612), .A2(n592), .ZN(n604) );
  NAND2_X1 U96 ( .A1(n622), .A2(n592), .ZN(n614) );
  NAND2_X1 U97 ( .A1(n672), .A2(n591), .ZN(n664) );
  NAND2_X1 U98 ( .A1(n672), .A2(n602), .ZN(n674) );
  NAND2_X1 U99 ( .A1(n672), .A2(n612), .ZN(n683) );
  NAND2_X1 U100 ( .A1(n672), .A2(n622), .ZN(n692) );
  NAND2_X1 U101 ( .A1(n745), .A2(n591), .ZN(n737) );
  NAND2_X1 U102 ( .A1(n745), .A2(n602), .ZN(n747) );
  NAND2_X1 U103 ( .A1(n745), .A2(n612), .ZN(n756) );
  NAND2_X1 U104 ( .A1(n745), .A2(n622), .ZN(n765) );
  NAND2_X1 U105 ( .A1(n818), .A2(n591), .ZN(n810) );
  NAND2_X1 U106 ( .A1(n818), .A2(n602), .ZN(n820) );
  NAND2_X1 U107 ( .A1(n818), .A2(n612), .ZN(n829) );
  NAND2_X1 U108 ( .A1(n818), .A2(n622), .ZN(n838) );
  NAND2_X1 U109 ( .A1(n891), .A2(n591), .ZN(n883) );
  NAND2_X1 U110 ( .A1(n891), .A2(n602), .ZN(n893) );
  NAND2_X1 U111 ( .A1(n891), .A2(n612), .ZN(n902) );
  NAND2_X1 U112 ( .A1(n891), .A2(n622), .ZN(n911) );
  NAND2_X1 U113 ( .A1(n964), .A2(n591), .ZN(n956) );
  NAND2_X1 U114 ( .A1(n964), .A2(n602), .ZN(n966) );
  NAND2_X1 U115 ( .A1(n964), .A2(n612), .ZN(n975) );
  NAND2_X1 U116 ( .A1(n964), .A2(n622), .ZN(n984) );
  NAND2_X1 U117 ( .A1(n1037), .A2(n591), .ZN(n1029) );
  NAND2_X1 U118 ( .A1(n1037), .A2(n602), .ZN(n1039) );
  NAND2_X1 U119 ( .A1(n1037), .A2(n612), .ZN(n1048) );
  NAND2_X1 U120 ( .A1(n1037), .A2(n622), .ZN(n1057) );
  NAND2_X1 U121 ( .A1(n1110), .A2(n591), .ZN(n1102) );
  NAND2_X1 U122 ( .A1(n1110), .A2(n602), .ZN(n1112) );
  NAND2_X1 U123 ( .A1(n1110), .A2(n612), .ZN(n1121) );
  NAND2_X1 U124 ( .A1(n1110), .A2(n622), .ZN(n1130) );
  NAND2_X1 U125 ( .A1(n672), .A2(n632), .ZN(n701) );
  NAND2_X1 U126 ( .A1(n672), .A2(n642), .ZN(n710) );
  NAND2_X1 U127 ( .A1(n672), .A2(n652), .ZN(n719) );
  NAND2_X1 U128 ( .A1(n672), .A2(n662), .ZN(n728) );
  NAND2_X1 U129 ( .A1(n745), .A2(n632), .ZN(n774) );
  NAND2_X1 U130 ( .A1(n745), .A2(n642), .ZN(n783) );
  NAND2_X1 U131 ( .A1(n745), .A2(n652), .ZN(n792) );
  NAND2_X1 U132 ( .A1(n745), .A2(n662), .ZN(n801) );
  NAND2_X1 U133 ( .A1(n818), .A2(n632), .ZN(n847) );
  NAND2_X1 U134 ( .A1(n818), .A2(n642), .ZN(n856) );
  NAND2_X1 U135 ( .A1(n818), .A2(n652), .ZN(n865) );
  NAND2_X1 U136 ( .A1(n818), .A2(n662), .ZN(n874) );
  NAND2_X1 U137 ( .A1(n891), .A2(n632), .ZN(n920) );
  NAND2_X1 U138 ( .A1(n891), .A2(n642), .ZN(n929) );
  NAND2_X1 U139 ( .A1(n891), .A2(n652), .ZN(n938) );
  NAND2_X1 U140 ( .A1(n891), .A2(n662), .ZN(n947) );
  NAND2_X1 U141 ( .A1(n964), .A2(n632), .ZN(n993) );
  NAND2_X1 U142 ( .A1(n964), .A2(n642), .ZN(n1002) );
  NAND2_X1 U143 ( .A1(n964), .A2(n652), .ZN(n1011) );
  NAND2_X1 U144 ( .A1(n964), .A2(n662), .ZN(n1020) );
  NAND2_X1 U145 ( .A1(n1037), .A2(n632), .ZN(n1066) );
  NAND2_X1 U146 ( .A1(n1037), .A2(n642), .ZN(n1075) );
  NAND2_X1 U147 ( .A1(n1037), .A2(n652), .ZN(n1084) );
  NAND2_X1 U148 ( .A1(n1037), .A2(n662), .ZN(n1093) );
  NAND2_X1 U149 ( .A1(n1110), .A2(n632), .ZN(n1139) );
  NAND2_X1 U150 ( .A1(n1110), .A2(n642), .ZN(n1148) );
  NAND2_X1 U151 ( .A1(n1110), .A2(n652), .ZN(n1157) );
  NAND2_X1 U152 ( .A1(n1110), .A2(n662), .ZN(n1166) );
  NAND2_X1 U153 ( .A1(n632), .A2(n592), .ZN(n624) );
  NAND2_X1 U154 ( .A1(n642), .A2(n592), .ZN(n634) );
  NAND2_X1 U155 ( .A1(n652), .A2(n592), .ZN(n644) );
  NAND2_X1 U156 ( .A1(n662), .A2(n592), .ZN(n654) );
  AND4_X1 U157 ( .A1(wr_en), .A2(n520), .A3(n521), .A4(n1690), .ZN(n592) );
  AND3_X1 U158 ( .A1(n518), .A2(n519), .A3(N12), .ZN(n632) );
  AND3_X1 U159 ( .A1(N11), .A2(n518), .A3(N12), .ZN(n652) );
  INV_X1 U160 ( .A(N15), .ZN(n1690) );
  INV_X1 U161 ( .A(n700), .ZN(n1529) );
  AOI22_X1 U162 ( .A1(data_in[0]), .A2(n1677), .B1(n701), .B2(\mem[12][0] ), 
        .ZN(n700) );
  INV_X1 U163 ( .A(n702), .ZN(n1528) );
  AOI22_X1 U164 ( .A1(data_in[1]), .A2(n1677), .B1(n701), .B2(\mem[12][1] ), 
        .ZN(n702) );
  INV_X1 U165 ( .A(n703), .ZN(n1527) );
  AOI22_X1 U166 ( .A1(data_in[2]), .A2(n1677), .B1(n701), .B2(\mem[12][2] ), 
        .ZN(n703) );
  INV_X1 U167 ( .A(n704), .ZN(n1526) );
  AOI22_X1 U168 ( .A1(data_in[3]), .A2(n1677), .B1(n701), .B2(\mem[12][3] ), 
        .ZN(n704) );
  INV_X1 U169 ( .A(n705), .ZN(n1525) );
  AOI22_X1 U170 ( .A1(data_in[4]), .A2(n1677), .B1(n701), .B2(\mem[12][4] ), 
        .ZN(n705) );
  INV_X1 U171 ( .A(n706), .ZN(n1524) );
  AOI22_X1 U172 ( .A1(data_in[5]), .A2(n1677), .B1(n701), .B2(\mem[12][5] ), 
        .ZN(n706) );
  INV_X1 U173 ( .A(n707), .ZN(n1523) );
  AOI22_X1 U174 ( .A1(data_in[6]), .A2(n1677), .B1(n701), .B2(\mem[12][6] ), 
        .ZN(n707) );
  INV_X1 U175 ( .A(n708), .ZN(n1522) );
  AOI22_X1 U176 ( .A1(data_in[7]), .A2(n1677), .B1(n701), .B2(\mem[12][7] ), 
        .ZN(n708) );
  INV_X1 U177 ( .A(n718), .ZN(n1513) );
  AOI22_X1 U178 ( .A1(data_in[0]), .A2(n1675), .B1(n719), .B2(\mem[14][0] ), 
        .ZN(n718) );
  INV_X1 U179 ( .A(n720), .ZN(n1512) );
  AOI22_X1 U180 ( .A1(data_in[1]), .A2(n1675), .B1(n719), .B2(\mem[14][1] ), 
        .ZN(n720) );
  INV_X1 U181 ( .A(n721), .ZN(n1511) );
  AOI22_X1 U182 ( .A1(data_in[2]), .A2(n1675), .B1(n719), .B2(\mem[14][2] ), 
        .ZN(n721) );
  INV_X1 U183 ( .A(n722), .ZN(n1510) );
  AOI22_X1 U184 ( .A1(data_in[3]), .A2(n1675), .B1(n719), .B2(\mem[14][3] ), 
        .ZN(n722) );
  INV_X1 U185 ( .A(n723), .ZN(n1509) );
  AOI22_X1 U186 ( .A1(data_in[4]), .A2(n1675), .B1(n719), .B2(\mem[14][4] ), 
        .ZN(n723) );
  INV_X1 U187 ( .A(n724), .ZN(n1508) );
  AOI22_X1 U188 ( .A1(data_in[5]), .A2(n1675), .B1(n719), .B2(\mem[14][5] ), 
        .ZN(n724) );
  INV_X1 U189 ( .A(n725), .ZN(n1507) );
  AOI22_X1 U190 ( .A1(data_in[6]), .A2(n1675), .B1(n719), .B2(\mem[14][6] ), 
        .ZN(n725) );
  INV_X1 U191 ( .A(n726), .ZN(n1506) );
  AOI22_X1 U192 ( .A1(data_in[7]), .A2(n1675), .B1(n719), .B2(\mem[14][7] ), 
        .ZN(n726) );
  INV_X1 U193 ( .A(n773), .ZN(n1465) );
  AOI22_X1 U194 ( .A1(data_in[0]), .A2(n1669), .B1(n774), .B2(\mem[20][0] ), 
        .ZN(n773) );
  INV_X1 U195 ( .A(n775), .ZN(n1464) );
  AOI22_X1 U196 ( .A1(data_in[1]), .A2(n1669), .B1(n774), .B2(\mem[20][1] ), 
        .ZN(n775) );
  INV_X1 U197 ( .A(n776), .ZN(n1463) );
  AOI22_X1 U198 ( .A1(data_in[2]), .A2(n1669), .B1(n774), .B2(\mem[20][2] ), 
        .ZN(n776) );
  INV_X1 U199 ( .A(n777), .ZN(n1462) );
  AOI22_X1 U200 ( .A1(data_in[3]), .A2(n1669), .B1(n774), .B2(\mem[20][3] ), 
        .ZN(n777) );
  INV_X1 U201 ( .A(n778), .ZN(n1461) );
  AOI22_X1 U202 ( .A1(data_in[4]), .A2(n1669), .B1(n774), .B2(\mem[20][4] ), 
        .ZN(n778) );
  INV_X1 U203 ( .A(n779), .ZN(n1460) );
  AOI22_X1 U204 ( .A1(data_in[5]), .A2(n1669), .B1(n774), .B2(\mem[20][5] ), 
        .ZN(n779) );
  INV_X1 U205 ( .A(n780), .ZN(n1459) );
  AOI22_X1 U206 ( .A1(data_in[6]), .A2(n1669), .B1(n774), .B2(\mem[20][6] ), 
        .ZN(n780) );
  INV_X1 U207 ( .A(n781), .ZN(n1458) );
  AOI22_X1 U208 ( .A1(data_in[7]), .A2(n1669), .B1(n774), .B2(\mem[20][7] ), 
        .ZN(n781) );
  INV_X1 U209 ( .A(n791), .ZN(n1449) );
  AOI22_X1 U210 ( .A1(data_in[0]), .A2(n1667), .B1(n792), .B2(\mem[22][0] ), 
        .ZN(n791) );
  INV_X1 U211 ( .A(n793), .ZN(n1448) );
  AOI22_X1 U212 ( .A1(data_in[1]), .A2(n1667), .B1(n792), .B2(\mem[22][1] ), 
        .ZN(n793) );
  INV_X1 U213 ( .A(n794), .ZN(n1447) );
  AOI22_X1 U214 ( .A1(data_in[2]), .A2(n1667), .B1(n792), .B2(\mem[22][2] ), 
        .ZN(n794) );
  INV_X1 U215 ( .A(n795), .ZN(n1446) );
  AOI22_X1 U216 ( .A1(data_in[3]), .A2(n1667), .B1(n792), .B2(\mem[22][3] ), 
        .ZN(n795) );
  INV_X1 U217 ( .A(n796), .ZN(n1445) );
  AOI22_X1 U218 ( .A1(data_in[4]), .A2(n1667), .B1(n792), .B2(\mem[22][4] ), 
        .ZN(n796) );
  INV_X1 U219 ( .A(n797), .ZN(n1444) );
  AOI22_X1 U220 ( .A1(data_in[5]), .A2(n1667), .B1(n792), .B2(\mem[22][5] ), 
        .ZN(n797) );
  INV_X1 U221 ( .A(n798), .ZN(n1443) );
  AOI22_X1 U222 ( .A1(data_in[6]), .A2(n1667), .B1(n792), .B2(\mem[22][6] ), 
        .ZN(n798) );
  INV_X1 U223 ( .A(n799), .ZN(n1442) );
  AOI22_X1 U224 ( .A1(data_in[7]), .A2(n1667), .B1(n792), .B2(\mem[22][7] ), 
        .ZN(n799) );
  INV_X1 U225 ( .A(n846), .ZN(n1401) );
  AOI22_X1 U226 ( .A1(data_in[0]), .A2(n1661), .B1(n847), .B2(\mem[28][0] ), 
        .ZN(n846) );
  INV_X1 U227 ( .A(n848), .ZN(n1400) );
  AOI22_X1 U228 ( .A1(data_in[1]), .A2(n1661), .B1(n847), .B2(\mem[28][1] ), 
        .ZN(n848) );
  INV_X1 U229 ( .A(n849), .ZN(n1399) );
  AOI22_X1 U230 ( .A1(data_in[2]), .A2(n1661), .B1(n847), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U231 ( .A(n850), .ZN(n1398) );
  AOI22_X1 U232 ( .A1(data_in[3]), .A2(n1661), .B1(n847), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U233 ( .A(n851), .ZN(n1397) );
  AOI22_X1 U234 ( .A1(data_in[4]), .A2(n1661), .B1(n847), .B2(\mem[28][4] ), 
        .ZN(n851) );
  INV_X1 U235 ( .A(n852), .ZN(n1396) );
  AOI22_X1 U236 ( .A1(data_in[5]), .A2(n1661), .B1(n847), .B2(\mem[28][5] ), 
        .ZN(n852) );
  INV_X1 U237 ( .A(n853), .ZN(n1395) );
  AOI22_X1 U238 ( .A1(data_in[6]), .A2(n1661), .B1(n847), .B2(\mem[28][6] ), 
        .ZN(n853) );
  INV_X1 U239 ( .A(n854), .ZN(n1394) );
  AOI22_X1 U240 ( .A1(data_in[7]), .A2(n1661), .B1(n847), .B2(\mem[28][7] ), 
        .ZN(n854) );
  INV_X1 U241 ( .A(n864), .ZN(n1385) );
  AOI22_X1 U242 ( .A1(data_in[0]), .A2(n1659), .B1(n865), .B2(\mem[30][0] ), 
        .ZN(n864) );
  INV_X1 U243 ( .A(n866), .ZN(n1384) );
  AOI22_X1 U244 ( .A1(data_in[1]), .A2(n1659), .B1(n865), .B2(\mem[30][1] ), 
        .ZN(n866) );
  INV_X1 U245 ( .A(n867), .ZN(n1383) );
  AOI22_X1 U246 ( .A1(data_in[2]), .A2(n1659), .B1(n865), .B2(\mem[30][2] ), 
        .ZN(n867) );
  INV_X1 U247 ( .A(n868), .ZN(n1382) );
  AOI22_X1 U248 ( .A1(data_in[3]), .A2(n1659), .B1(n865), .B2(\mem[30][3] ), 
        .ZN(n868) );
  INV_X1 U249 ( .A(n869), .ZN(n1381) );
  AOI22_X1 U250 ( .A1(data_in[4]), .A2(n1659), .B1(n865), .B2(\mem[30][4] ), 
        .ZN(n869) );
  INV_X1 U251 ( .A(n870), .ZN(n1380) );
  AOI22_X1 U252 ( .A1(data_in[5]), .A2(n1659), .B1(n865), .B2(\mem[30][5] ), 
        .ZN(n870) );
  INV_X1 U253 ( .A(n871), .ZN(n1379) );
  AOI22_X1 U254 ( .A1(data_in[6]), .A2(n1659), .B1(n865), .B2(\mem[30][6] ), 
        .ZN(n871) );
  INV_X1 U255 ( .A(n872), .ZN(n1378) );
  AOI22_X1 U256 ( .A1(data_in[7]), .A2(n1659), .B1(n865), .B2(\mem[30][7] ), 
        .ZN(n872) );
  INV_X1 U257 ( .A(n919), .ZN(n1337) );
  AOI22_X1 U258 ( .A1(data_in[0]), .A2(n1653), .B1(n920), .B2(\mem[36][0] ), 
        .ZN(n919) );
  INV_X1 U259 ( .A(n921), .ZN(n1336) );
  AOI22_X1 U260 ( .A1(data_in[1]), .A2(n1653), .B1(n920), .B2(\mem[36][1] ), 
        .ZN(n921) );
  INV_X1 U261 ( .A(n922), .ZN(n1335) );
  AOI22_X1 U262 ( .A1(data_in[2]), .A2(n1653), .B1(n920), .B2(\mem[36][2] ), 
        .ZN(n922) );
  INV_X1 U263 ( .A(n923), .ZN(n1334) );
  AOI22_X1 U264 ( .A1(data_in[3]), .A2(n1653), .B1(n920), .B2(\mem[36][3] ), 
        .ZN(n923) );
  INV_X1 U265 ( .A(n924), .ZN(n1333) );
  AOI22_X1 U266 ( .A1(data_in[4]), .A2(n1653), .B1(n920), .B2(\mem[36][4] ), 
        .ZN(n924) );
  INV_X1 U267 ( .A(n925), .ZN(n1332) );
  AOI22_X1 U268 ( .A1(data_in[5]), .A2(n1653), .B1(n920), .B2(\mem[36][5] ), 
        .ZN(n925) );
  INV_X1 U269 ( .A(n926), .ZN(n1331) );
  AOI22_X1 U270 ( .A1(data_in[6]), .A2(n1653), .B1(n920), .B2(\mem[36][6] ), 
        .ZN(n926) );
  INV_X1 U271 ( .A(n927), .ZN(n1330) );
  AOI22_X1 U272 ( .A1(data_in[7]), .A2(n1653), .B1(n920), .B2(\mem[36][7] ), 
        .ZN(n927) );
  INV_X1 U273 ( .A(n937), .ZN(n1321) );
  AOI22_X1 U274 ( .A1(data_in[0]), .A2(n1651), .B1(n938), .B2(\mem[38][0] ), 
        .ZN(n937) );
  INV_X1 U275 ( .A(n939), .ZN(n1320) );
  AOI22_X1 U276 ( .A1(data_in[1]), .A2(n1651), .B1(n938), .B2(\mem[38][1] ), 
        .ZN(n939) );
  INV_X1 U277 ( .A(n940), .ZN(n1319) );
  AOI22_X1 U278 ( .A1(data_in[2]), .A2(n1651), .B1(n938), .B2(\mem[38][2] ), 
        .ZN(n940) );
  INV_X1 U279 ( .A(n941), .ZN(n1318) );
  AOI22_X1 U280 ( .A1(data_in[3]), .A2(n1651), .B1(n938), .B2(\mem[38][3] ), 
        .ZN(n941) );
  INV_X1 U281 ( .A(n942), .ZN(n1317) );
  AOI22_X1 U282 ( .A1(data_in[4]), .A2(n1651), .B1(n938), .B2(\mem[38][4] ), 
        .ZN(n942) );
  INV_X1 U283 ( .A(n943), .ZN(n1316) );
  AOI22_X1 U284 ( .A1(data_in[5]), .A2(n1651), .B1(n938), .B2(\mem[38][5] ), 
        .ZN(n943) );
  INV_X1 U285 ( .A(n944), .ZN(n1315) );
  AOI22_X1 U286 ( .A1(data_in[6]), .A2(n1651), .B1(n938), .B2(\mem[38][6] ), 
        .ZN(n944) );
  INV_X1 U287 ( .A(n945), .ZN(n1314) );
  AOI22_X1 U288 ( .A1(data_in[7]), .A2(n1651), .B1(n938), .B2(\mem[38][7] ), 
        .ZN(n945) );
  INV_X1 U289 ( .A(n992), .ZN(n1273) );
  AOI22_X1 U290 ( .A1(data_in[0]), .A2(n1645), .B1(n993), .B2(\mem[44][0] ), 
        .ZN(n992) );
  INV_X1 U291 ( .A(n994), .ZN(n1272) );
  AOI22_X1 U292 ( .A1(data_in[1]), .A2(n1645), .B1(n993), .B2(\mem[44][1] ), 
        .ZN(n994) );
  INV_X1 U293 ( .A(n995), .ZN(n1271) );
  AOI22_X1 U294 ( .A1(data_in[2]), .A2(n1645), .B1(n993), .B2(\mem[44][2] ), 
        .ZN(n995) );
  INV_X1 U295 ( .A(n996), .ZN(n1270) );
  AOI22_X1 U296 ( .A1(data_in[3]), .A2(n1645), .B1(n993), .B2(\mem[44][3] ), 
        .ZN(n996) );
  INV_X1 U297 ( .A(n997), .ZN(n1269) );
  AOI22_X1 U298 ( .A1(data_in[4]), .A2(n1645), .B1(n993), .B2(\mem[44][4] ), 
        .ZN(n997) );
  INV_X1 U299 ( .A(n998), .ZN(n1268) );
  AOI22_X1 U300 ( .A1(data_in[5]), .A2(n1645), .B1(n993), .B2(\mem[44][5] ), 
        .ZN(n998) );
  INV_X1 U301 ( .A(n999), .ZN(n1267) );
  AOI22_X1 U302 ( .A1(data_in[6]), .A2(n1645), .B1(n993), .B2(\mem[44][6] ), 
        .ZN(n999) );
  INV_X1 U303 ( .A(n1000), .ZN(n1266) );
  AOI22_X1 U304 ( .A1(data_in[7]), .A2(n1645), .B1(n993), .B2(\mem[44][7] ), 
        .ZN(n1000) );
  INV_X1 U305 ( .A(n1010), .ZN(n1257) );
  AOI22_X1 U306 ( .A1(data_in[0]), .A2(n1643), .B1(n1011), .B2(\mem[46][0] ), 
        .ZN(n1010) );
  INV_X1 U307 ( .A(n1012), .ZN(n1256) );
  AOI22_X1 U308 ( .A1(data_in[1]), .A2(n1643), .B1(n1011), .B2(\mem[46][1] ), 
        .ZN(n1012) );
  INV_X1 U309 ( .A(n1013), .ZN(n1255) );
  AOI22_X1 U310 ( .A1(data_in[2]), .A2(n1643), .B1(n1011), .B2(\mem[46][2] ), 
        .ZN(n1013) );
  INV_X1 U311 ( .A(n1014), .ZN(n1254) );
  AOI22_X1 U312 ( .A1(data_in[3]), .A2(n1643), .B1(n1011), .B2(\mem[46][3] ), 
        .ZN(n1014) );
  INV_X1 U313 ( .A(n1015), .ZN(n1253) );
  AOI22_X1 U314 ( .A1(data_in[4]), .A2(n1643), .B1(n1011), .B2(\mem[46][4] ), 
        .ZN(n1015) );
  INV_X1 U315 ( .A(n1016), .ZN(n1252) );
  AOI22_X1 U316 ( .A1(data_in[5]), .A2(n1643), .B1(n1011), .B2(\mem[46][5] ), 
        .ZN(n1016) );
  INV_X1 U317 ( .A(n1017), .ZN(n1251) );
  AOI22_X1 U318 ( .A1(data_in[6]), .A2(n1643), .B1(n1011), .B2(\mem[46][6] ), 
        .ZN(n1017) );
  INV_X1 U319 ( .A(n1018), .ZN(n1250) );
  AOI22_X1 U320 ( .A1(data_in[7]), .A2(n1643), .B1(n1011), .B2(\mem[46][7] ), 
        .ZN(n1018) );
  INV_X1 U321 ( .A(n1065), .ZN(n1209) );
  AOI22_X1 U322 ( .A1(data_in[0]), .A2(n1637), .B1(n1066), .B2(\mem[52][0] ), 
        .ZN(n1065) );
  INV_X1 U323 ( .A(n1067), .ZN(n1208) );
  AOI22_X1 U324 ( .A1(data_in[1]), .A2(n1637), .B1(n1066), .B2(\mem[52][1] ), 
        .ZN(n1067) );
  INV_X1 U325 ( .A(n1068), .ZN(n1207) );
  AOI22_X1 U326 ( .A1(data_in[2]), .A2(n1637), .B1(n1066), .B2(\mem[52][2] ), 
        .ZN(n1068) );
  INV_X1 U327 ( .A(n1069), .ZN(n1206) );
  AOI22_X1 U328 ( .A1(data_in[3]), .A2(n1637), .B1(n1066), .B2(\mem[52][3] ), 
        .ZN(n1069) );
  INV_X1 U329 ( .A(n1070), .ZN(n1205) );
  AOI22_X1 U330 ( .A1(data_in[4]), .A2(n1637), .B1(n1066), .B2(\mem[52][4] ), 
        .ZN(n1070) );
  INV_X1 U331 ( .A(n1071), .ZN(n1204) );
  AOI22_X1 U332 ( .A1(data_in[5]), .A2(n1637), .B1(n1066), .B2(\mem[52][5] ), 
        .ZN(n1071) );
  INV_X1 U333 ( .A(n1072), .ZN(n1203) );
  AOI22_X1 U334 ( .A1(data_in[6]), .A2(n1637), .B1(n1066), .B2(\mem[52][6] ), 
        .ZN(n1072) );
  INV_X1 U335 ( .A(n1073), .ZN(n1202) );
  AOI22_X1 U336 ( .A1(data_in[7]), .A2(n1637), .B1(n1066), .B2(\mem[52][7] ), 
        .ZN(n1073) );
  INV_X1 U337 ( .A(n1083), .ZN(n1193) );
  AOI22_X1 U338 ( .A1(data_in[0]), .A2(n1635), .B1(n1084), .B2(\mem[54][0] ), 
        .ZN(n1083) );
  INV_X1 U339 ( .A(n1085), .ZN(n1192) );
  AOI22_X1 U340 ( .A1(data_in[1]), .A2(n1635), .B1(n1084), .B2(\mem[54][1] ), 
        .ZN(n1085) );
  INV_X1 U341 ( .A(n1086), .ZN(n1191) );
  AOI22_X1 U342 ( .A1(data_in[2]), .A2(n1635), .B1(n1084), .B2(\mem[54][2] ), 
        .ZN(n1086) );
  INV_X1 U343 ( .A(n1087), .ZN(n1190) );
  AOI22_X1 U344 ( .A1(data_in[3]), .A2(n1635), .B1(n1084), .B2(\mem[54][3] ), 
        .ZN(n1087) );
  INV_X1 U345 ( .A(n1088), .ZN(n1189) );
  AOI22_X1 U346 ( .A1(data_in[4]), .A2(n1635), .B1(n1084), .B2(\mem[54][4] ), 
        .ZN(n1088) );
  INV_X1 U347 ( .A(n1089), .ZN(n1188) );
  AOI22_X1 U348 ( .A1(data_in[5]), .A2(n1635), .B1(n1084), .B2(\mem[54][5] ), 
        .ZN(n1089) );
  INV_X1 U349 ( .A(n1090), .ZN(n1187) );
  AOI22_X1 U350 ( .A1(data_in[6]), .A2(n1635), .B1(n1084), .B2(\mem[54][6] ), 
        .ZN(n1090) );
  INV_X1 U351 ( .A(n1091), .ZN(n1186) );
  AOI22_X1 U352 ( .A1(data_in[7]), .A2(n1635), .B1(n1084), .B2(\mem[54][7] ), 
        .ZN(n1091) );
  INV_X1 U353 ( .A(n1138), .ZN(n553) );
  AOI22_X1 U354 ( .A1(data_in[0]), .A2(n1629), .B1(n1139), .B2(\mem[60][0] ), 
        .ZN(n1138) );
  INV_X1 U355 ( .A(n1140), .ZN(n552) );
  AOI22_X1 U356 ( .A1(data_in[1]), .A2(n1629), .B1(n1139), .B2(\mem[60][1] ), 
        .ZN(n1140) );
  INV_X1 U357 ( .A(n1141), .ZN(n551) );
  AOI22_X1 U358 ( .A1(data_in[2]), .A2(n1629), .B1(n1139), .B2(\mem[60][2] ), 
        .ZN(n1141) );
  INV_X1 U359 ( .A(n1142), .ZN(n550) );
  AOI22_X1 U360 ( .A1(data_in[3]), .A2(n1629), .B1(n1139), .B2(\mem[60][3] ), 
        .ZN(n1142) );
  INV_X1 U361 ( .A(n1143), .ZN(n549) );
  AOI22_X1 U362 ( .A1(data_in[4]), .A2(n1629), .B1(n1139), .B2(\mem[60][4] ), 
        .ZN(n1143) );
  INV_X1 U363 ( .A(n1144), .ZN(n548) );
  AOI22_X1 U364 ( .A1(data_in[5]), .A2(n1629), .B1(n1139), .B2(\mem[60][5] ), 
        .ZN(n1144) );
  INV_X1 U365 ( .A(n1145), .ZN(n547) );
  AOI22_X1 U366 ( .A1(data_in[6]), .A2(n1629), .B1(n1139), .B2(\mem[60][6] ), 
        .ZN(n1145) );
  INV_X1 U367 ( .A(n1146), .ZN(n546) );
  AOI22_X1 U368 ( .A1(data_in[7]), .A2(n1629), .B1(n1139), .B2(\mem[60][7] ), 
        .ZN(n1146) );
  INV_X1 U369 ( .A(n1156), .ZN(n537) );
  AOI22_X1 U370 ( .A1(data_in[0]), .A2(n1627), .B1(n1157), .B2(\mem[62][0] ), 
        .ZN(n1156) );
  INV_X1 U371 ( .A(n1158), .ZN(n536) );
  AOI22_X1 U372 ( .A1(data_in[1]), .A2(n1627), .B1(n1157), .B2(\mem[62][1] ), 
        .ZN(n1158) );
  INV_X1 U373 ( .A(n1159), .ZN(n535) );
  AOI22_X1 U374 ( .A1(data_in[2]), .A2(n1627), .B1(n1157), .B2(\mem[62][2] ), 
        .ZN(n1159) );
  INV_X1 U375 ( .A(n1160), .ZN(n534) );
  AOI22_X1 U376 ( .A1(data_in[3]), .A2(n1627), .B1(n1157), .B2(\mem[62][3] ), 
        .ZN(n1160) );
  INV_X1 U377 ( .A(n1161), .ZN(n533) );
  AOI22_X1 U378 ( .A1(data_in[4]), .A2(n1627), .B1(n1157), .B2(\mem[62][4] ), 
        .ZN(n1161) );
  INV_X1 U379 ( .A(n1162), .ZN(n532) );
  AOI22_X1 U380 ( .A1(data_in[5]), .A2(n1627), .B1(n1157), .B2(\mem[62][5] ), 
        .ZN(n1162) );
  INV_X1 U381 ( .A(n1163), .ZN(n531) );
  AOI22_X1 U382 ( .A1(data_in[6]), .A2(n1627), .B1(n1157), .B2(\mem[62][6] ), 
        .ZN(n1163) );
  INV_X1 U383 ( .A(n1164), .ZN(n530) );
  AOI22_X1 U384 ( .A1(data_in[7]), .A2(n1627), .B1(n1157), .B2(\mem[62][7] ), 
        .ZN(n1164) );
  INV_X1 U385 ( .A(N14), .ZN(n521) );
  INV_X1 U386 ( .A(N13), .ZN(n520) );
  INV_X1 U387 ( .A(n663), .ZN(n1561) );
  AOI22_X1 U388 ( .A1(data_in[0]), .A2(n1681), .B1(n664), .B2(\mem[8][0] ), 
        .ZN(n663) );
  INV_X1 U389 ( .A(n665), .ZN(n1560) );
  AOI22_X1 U390 ( .A1(data_in[1]), .A2(n1681), .B1(n664), .B2(\mem[8][1] ), 
        .ZN(n665) );
  INV_X1 U391 ( .A(n666), .ZN(n1559) );
  AOI22_X1 U392 ( .A1(data_in[2]), .A2(n1681), .B1(n664), .B2(\mem[8][2] ), 
        .ZN(n666) );
  INV_X1 U393 ( .A(n667), .ZN(n1558) );
  AOI22_X1 U394 ( .A1(data_in[3]), .A2(n1681), .B1(n664), .B2(\mem[8][3] ), 
        .ZN(n667) );
  INV_X1 U395 ( .A(n668), .ZN(n1557) );
  AOI22_X1 U396 ( .A1(data_in[4]), .A2(n1681), .B1(n664), .B2(\mem[8][4] ), 
        .ZN(n668) );
  INV_X1 U397 ( .A(n669), .ZN(n1556) );
  AOI22_X1 U398 ( .A1(data_in[5]), .A2(n1681), .B1(n664), .B2(\mem[8][5] ), 
        .ZN(n669) );
  INV_X1 U399 ( .A(n670), .ZN(n1555) );
  AOI22_X1 U400 ( .A1(data_in[6]), .A2(n1681), .B1(n664), .B2(\mem[8][6] ), 
        .ZN(n670) );
  INV_X1 U401 ( .A(n671), .ZN(n1554) );
  AOI22_X1 U402 ( .A1(data_in[7]), .A2(n1681), .B1(n664), .B2(\mem[8][7] ), 
        .ZN(n671) );
  INV_X1 U403 ( .A(n673), .ZN(n1553) );
  AOI22_X1 U404 ( .A1(data_in[0]), .A2(n1680), .B1(n674), .B2(\mem[9][0] ), 
        .ZN(n673) );
  INV_X1 U405 ( .A(n675), .ZN(n1552) );
  AOI22_X1 U406 ( .A1(data_in[1]), .A2(n1680), .B1(n674), .B2(\mem[9][1] ), 
        .ZN(n675) );
  INV_X1 U407 ( .A(n676), .ZN(n1551) );
  AOI22_X1 U408 ( .A1(data_in[2]), .A2(n1680), .B1(n674), .B2(\mem[9][2] ), 
        .ZN(n676) );
  INV_X1 U409 ( .A(n677), .ZN(n1550) );
  AOI22_X1 U410 ( .A1(data_in[3]), .A2(n1680), .B1(n674), .B2(\mem[9][3] ), 
        .ZN(n677) );
  INV_X1 U411 ( .A(n678), .ZN(n1549) );
  AOI22_X1 U412 ( .A1(data_in[4]), .A2(n1680), .B1(n674), .B2(\mem[9][4] ), 
        .ZN(n678) );
  INV_X1 U413 ( .A(n679), .ZN(n1548) );
  AOI22_X1 U414 ( .A1(data_in[5]), .A2(n1680), .B1(n674), .B2(\mem[9][5] ), 
        .ZN(n679) );
  INV_X1 U415 ( .A(n680), .ZN(n1547) );
  AOI22_X1 U416 ( .A1(data_in[6]), .A2(n1680), .B1(n674), .B2(\mem[9][6] ), 
        .ZN(n680) );
  INV_X1 U417 ( .A(n681), .ZN(n1546) );
  AOI22_X1 U418 ( .A1(data_in[7]), .A2(n1680), .B1(n674), .B2(\mem[9][7] ), 
        .ZN(n681) );
  INV_X1 U419 ( .A(n682), .ZN(n1545) );
  AOI22_X1 U420 ( .A1(data_in[0]), .A2(n1679), .B1(n683), .B2(\mem[10][0] ), 
        .ZN(n682) );
  INV_X1 U421 ( .A(n684), .ZN(n1544) );
  AOI22_X1 U422 ( .A1(data_in[1]), .A2(n1679), .B1(n683), .B2(\mem[10][1] ), 
        .ZN(n684) );
  INV_X1 U423 ( .A(n685), .ZN(n1543) );
  AOI22_X1 U424 ( .A1(data_in[2]), .A2(n1679), .B1(n683), .B2(\mem[10][2] ), 
        .ZN(n685) );
  INV_X1 U425 ( .A(n686), .ZN(n1542) );
  AOI22_X1 U426 ( .A1(data_in[3]), .A2(n1679), .B1(n683), .B2(\mem[10][3] ), 
        .ZN(n686) );
  INV_X1 U427 ( .A(n687), .ZN(n1541) );
  AOI22_X1 U428 ( .A1(data_in[4]), .A2(n1679), .B1(n683), .B2(\mem[10][4] ), 
        .ZN(n687) );
  INV_X1 U429 ( .A(n688), .ZN(n1540) );
  AOI22_X1 U430 ( .A1(data_in[5]), .A2(n1679), .B1(n683), .B2(\mem[10][5] ), 
        .ZN(n688) );
  INV_X1 U431 ( .A(n689), .ZN(n1539) );
  AOI22_X1 U432 ( .A1(data_in[6]), .A2(n1679), .B1(n683), .B2(\mem[10][6] ), 
        .ZN(n689) );
  INV_X1 U433 ( .A(n690), .ZN(n1538) );
  AOI22_X1 U434 ( .A1(data_in[7]), .A2(n1679), .B1(n683), .B2(\mem[10][7] ), 
        .ZN(n690) );
  INV_X1 U435 ( .A(n691), .ZN(n1537) );
  AOI22_X1 U436 ( .A1(data_in[0]), .A2(n1678), .B1(n692), .B2(\mem[11][0] ), 
        .ZN(n691) );
  INV_X1 U437 ( .A(n693), .ZN(n1536) );
  AOI22_X1 U438 ( .A1(data_in[1]), .A2(n1678), .B1(n692), .B2(\mem[11][1] ), 
        .ZN(n693) );
  INV_X1 U439 ( .A(n694), .ZN(n1535) );
  AOI22_X1 U440 ( .A1(data_in[2]), .A2(n1678), .B1(n692), .B2(\mem[11][2] ), 
        .ZN(n694) );
  INV_X1 U441 ( .A(n695), .ZN(n1534) );
  AOI22_X1 U442 ( .A1(data_in[3]), .A2(n1678), .B1(n692), .B2(\mem[11][3] ), 
        .ZN(n695) );
  INV_X1 U443 ( .A(n696), .ZN(n1533) );
  AOI22_X1 U444 ( .A1(data_in[4]), .A2(n1678), .B1(n692), .B2(\mem[11][4] ), 
        .ZN(n696) );
  INV_X1 U445 ( .A(n697), .ZN(n1532) );
  AOI22_X1 U446 ( .A1(data_in[5]), .A2(n1678), .B1(n692), .B2(\mem[11][5] ), 
        .ZN(n697) );
  INV_X1 U447 ( .A(n698), .ZN(n1531) );
  AOI22_X1 U448 ( .A1(data_in[6]), .A2(n1678), .B1(n692), .B2(\mem[11][6] ), 
        .ZN(n698) );
  INV_X1 U449 ( .A(n699), .ZN(n1530) );
  AOI22_X1 U450 ( .A1(data_in[7]), .A2(n1678), .B1(n692), .B2(\mem[11][7] ), 
        .ZN(n699) );
  INV_X1 U451 ( .A(n736), .ZN(n1497) );
  AOI22_X1 U452 ( .A1(data_in[0]), .A2(n1673), .B1(n737), .B2(\mem[16][0] ), 
        .ZN(n736) );
  INV_X1 U453 ( .A(n738), .ZN(n1496) );
  AOI22_X1 U454 ( .A1(data_in[1]), .A2(n1673), .B1(n737), .B2(\mem[16][1] ), 
        .ZN(n738) );
  INV_X1 U455 ( .A(n739), .ZN(n1495) );
  AOI22_X1 U456 ( .A1(data_in[2]), .A2(n1673), .B1(n737), .B2(\mem[16][2] ), 
        .ZN(n739) );
  INV_X1 U457 ( .A(n740), .ZN(n1494) );
  AOI22_X1 U458 ( .A1(data_in[3]), .A2(n1673), .B1(n737), .B2(\mem[16][3] ), 
        .ZN(n740) );
  INV_X1 U459 ( .A(n741), .ZN(n1493) );
  AOI22_X1 U460 ( .A1(data_in[4]), .A2(n1673), .B1(n737), .B2(\mem[16][4] ), 
        .ZN(n741) );
  INV_X1 U461 ( .A(n742), .ZN(n1492) );
  AOI22_X1 U462 ( .A1(data_in[5]), .A2(n1673), .B1(n737), .B2(\mem[16][5] ), 
        .ZN(n742) );
  INV_X1 U463 ( .A(n743), .ZN(n1491) );
  AOI22_X1 U464 ( .A1(data_in[6]), .A2(n1673), .B1(n737), .B2(\mem[16][6] ), 
        .ZN(n743) );
  INV_X1 U465 ( .A(n744), .ZN(n1490) );
  AOI22_X1 U466 ( .A1(data_in[7]), .A2(n1673), .B1(n737), .B2(\mem[16][7] ), 
        .ZN(n744) );
  INV_X1 U467 ( .A(n746), .ZN(n1489) );
  AOI22_X1 U468 ( .A1(data_in[0]), .A2(n1672), .B1(n747), .B2(\mem[17][0] ), 
        .ZN(n746) );
  INV_X1 U469 ( .A(n748), .ZN(n1488) );
  AOI22_X1 U470 ( .A1(data_in[1]), .A2(n1672), .B1(n747), .B2(\mem[17][1] ), 
        .ZN(n748) );
  INV_X1 U471 ( .A(n749), .ZN(n1487) );
  AOI22_X1 U472 ( .A1(data_in[2]), .A2(n1672), .B1(n747), .B2(\mem[17][2] ), 
        .ZN(n749) );
  INV_X1 U473 ( .A(n750), .ZN(n1486) );
  AOI22_X1 U474 ( .A1(data_in[3]), .A2(n1672), .B1(n747), .B2(\mem[17][3] ), 
        .ZN(n750) );
  INV_X1 U475 ( .A(n751), .ZN(n1485) );
  AOI22_X1 U476 ( .A1(data_in[4]), .A2(n1672), .B1(n747), .B2(\mem[17][4] ), 
        .ZN(n751) );
  INV_X1 U477 ( .A(n752), .ZN(n1484) );
  AOI22_X1 U478 ( .A1(data_in[5]), .A2(n1672), .B1(n747), .B2(\mem[17][5] ), 
        .ZN(n752) );
  INV_X1 U479 ( .A(n753), .ZN(n1483) );
  AOI22_X1 U480 ( .A1(data_in[6]), .A2(n1672), .B1(n747), .B2(\mem[17][6] ), 
        .ZN(n753) );
  INV_X1 U481 ( .A(n754), .ZN(n1482) );
  AOI22_X1 U482 ( .A1(data_in[7]), .A2(n1672), .B1(n747), .B2(\mem[17][7] ), 
        .ZN(n754) );
  INV_X1 U483 ( .A(n755), .ZN(n1481) );
  AOI22_X1 U484 ( .A1(data_in[0]), .A2(n1671), .B1(n756), .B2(\mem[18][0] ), 
        .ZN(n755) );
  INV_X1 U485 ( .A(n757), .ZN(n1480) );
  AOI22_X1 U486 ( .A1(data_in[1]), .A2(n1671), .B1(n756), .B2(\mem[18][1] ), 
        .ZN(n757) );
  INV_X1 U487 ( .A(n758), .ZN(n1479) );
  AOI22_X1 U488 ( .A1(data_in[2]), .A2(n1671), .B1(n756), .B2(\mem[18][2] ), 
        .ZN(n758) );
  INV_X1 U489 ( .A(n759), .ZN(n1478) );
  AOI22_X1 U490 ( .A1(data_in[3]), .A2(n1671), .B1(n756), .B2(\mem[18][3] ), 
        .ZN(n759) );
  INV_X1 U491 ( .A(n760), .ZN(n1477) );
  AOI22_X1 U492 ( .A1(data_in[4]), .A2(n1671), .B1(n756), .B2(\mem[18][4] ), 
        .ZN(n760) );
  INV_X1 U493 ( .A(n761), .ZN(n1476) );
  AOI22_X1 U494 ( .A1(data_in[5]), .A2(n1671), .B1(n756), .B2(\mem[18][5] ), 
        .ZN(n761) );
  INV_X1 U495 ( .A(n762), .ZN(n1475) );
  AOI22_X1 U496 ( .A1(data_in[6]), .A2(n1671), .B1(n756), .B2(\mem[18][6] ), 
        .ZN(n762) );
  INV_X1 U497 ( .A(n763), .ZN(n1474) );
  AOI22_X1 U498 ( .A1(data_in[7]), .A2(n1671), .B1(n756), .B2(\mem[18][7] ), 
        .ZN(n763) );
  INV_X1 U499 ( .A(n764), .ZN(n1473) );
  AOI22_X1 U500 ( .A1(data_in[0]), .A2(n1670), .B1(n765), .B2(\mem[19][0] ), 
        .ZN(n764) );
  INV_X1 U501 ( .A(n766), .ZN(n1472) );
  AOI22_X1 U502 ( .A1(data_in[1]), .A2(n1670), .B1(n765), .B2(\mem[19][1] ), 
        .ZN(n766) );
  INV_X1 U503 ( .A(n767), .ZN(n1471) );
  AOI22_X1 U504 ( .A1(data_in[2]), .A2(n1670), .B1(n765), .B2(\mem[19][2] ), 
        .ZN(n767) );
  INV_X1 U505 ( .A(n768), .ZN(n1470) );
  AOI22_X1 U506 ( .A1(data_in[3]), .A2(n1670), .B1(n765), .B2(\mem[19][3] ), 
        .ZN(n768) );
  INV_X1 U507 ( .A(n769), .ZN(n1469) );
  AOI22_X1 U508 ( .A1(data_in[4]), .A2(n1670), .B1(n765), .B2(\mem[19][4] ), 
        .ZN(n769) );
  INV_X1 U509 ( .A(n770), .ZN(n1468) );
  AOI22_X1 U510 ( .A1(data_in[5]), .A2(n1670), .B1(n765), .B2(\mem[19][5] ), 
        .ZN(n770) );
  INV_X1 U511 ( .A(n771), .ZN(n1467) );
  AOI22_X1 U512 ( .A1(data_in[6]), .A2(n1670), .B1(n765), .B2(\mem[19][6] ), 
        .ZN(n771) );
  INV_X1 U513 ( .A(n772), .ZN(n1466) );
  AOI22_X1 U514 ( .A1(data_in[7]), .A2(n1670), .B1(n765), .B2(\mem[19][7] ), 
        .ZN(n772) );
  INV_X1 U515 ( .A(n809), .ZN(n1433) );
  AOI22_X1 U516 ( .A1(data_in[0]), .A2(n1665), .B1(n810), .B2(\mem[24][0] ), 
        .ZN(n809) );
  INV_X1 U517 ( .A(n811), .ZN(n1432) );
  AOI22_X1 U518 ( .A1(data_in[1]), .A2(n1665), .B1(n810), .B2(\mem[24][1] ), 
        .ZN(n811) );
  INV_X1 U519 ( .A(n812), .ZN(n1431) );
  AOI22_X1 U520 ( .A1(data_in[2]), .A2(n1665), .B1(n810), .B2(\mem[24][2] ), 
        .ZN(n812) );
  INV_X1 U521 ( .A(n813), .ZN(n1430) );
  AOI22_X1 U522 ( .A1(data_in[3]), .A2(n1665), .B1(n810), .B2(\mem[24][3] ), 
        .ZN(n813) );
  INV_X1 U524 ( .A(n814), .ZN(n1429) );
  AOI22_X1 U525 ( .A1(data_in[4]), .A2(n1665), .B1(n810), .B2(\mem[24][4] ), 
        .ZN(n814) );
  INV_X1 U526 ( .A(n815), .ZN(n1428) );
  AOI22_X1 U527 ( .A1(data_in[5]), .A2(n1665), .B1(n810), .B2(\mem[24][5] ), 
        .ZN(n815) );
  INV_X1 U528 ( .A(n816), .ZN(n1427) );
  AOI22_X1 U529 ( .A1(data_in[6]), .A2(n1665), .B1(n810), .B2(\mem[24][6] ), 
        .ZN(n816) );
  INV_X1 U530 ( .A(n817), .ZN(n1426) );
  AOI22_X1 U531 ( .A1(data_in[7]), .A2(n1665), .B1(n810), .B2(\mem[24][7] ), 
        .ZN(n817) );
  INV_X1 U532 ( .A(n819), .ZN(n1425) );
  AOI22_X1 U534 ( .A1(data_in[0]), .A2(n1664), .B1(n820), .B2(\mem[25][0] ), 
        .ZN(n819) );
  INV_X1 U535 ( .A(n821), .ZN(n1424) );
  AOI22_X1 U536 ( .A1(data_in[1]), .A2(n1664), .B1(n820), .B2(\mem[25][1] ), 
        .ZN(n821) );
  INV_X1 U537 ( .A(n822), .ZN(n1423) );
  AOI22_X1 U538 ( .A1(data_in[2]), .A2(n1664), .B1(n820), .B2(\mem[25][2] ), 
        .ZN(n822) );
  INV_X1 U539 ( .A(n823), .ZN(n1422) );
  AOI22_X1 U540 ( .A1(data_in[3]), .A2(n1664), .B1(n820), .B2(\mem[25][3] ), 
        .ZN(n823) );
  INV_X1 U541 ( .A(n824), .ZN(n1421) );
  AOI22_X1 U542 ( .A1(data_in[4]), .A2(n1664), .B1(n820), .B2(\mem[25][4] ), 
        .ZN(n824) );
  INV_X1 U544 ( .A(n825), .ZN(n1420) );
  AOI22_X1 U545 ( .A1(data_in[5]), .A2(n1664), .B1(n820), .B2(\mem[25][5] ), 
        .ZN(n825) );
  INV_X1 U546 ( .A(n826), .ZN(n1419) );
  AOI22_X1 U547 ( .A1(data_in[6]), .A2(n1664), .B1(n820), .B2(\mem[25][6] ), 
        .ZN(n826) );
  INV_X1 U548 ( .A(n827), .ZN(n1418) );
  AOI22_X1 U549 ( .A1(data_in[7]), .A2(n1664), .B1(n820), .B2(\mem[25][7] ), 
        .ZN(n827) );
  INV_X1 U550 ( .A(n828), .ZN(n1417) );
  AOI22_X1 U551 ( .A1(data_in[0]), .A2(n1663), .B1(n829), .B2(\mem[26][0] ), 
        .ZN(n828) );
  INV_X1 U552 ( .A(n830), .ZN(n1416) );
  AOI22_X1 U554 ( .A1(data_in[1]), .A2(n1663), .B1(n829), .B2(\mem[26][1] ), 
        .ZN(n830) );
  INV_X1 U555 ( .A(n831), .ZN(n1415) );
  AOI22_X1 U556 ( .A1(data_in[2]), .A2(n1663), .B1(n829), .B2(\mem[26][2] ), 
        .ZN(n831) );
  INV_X1 U557 ( .A(n832), .ZN(n1414) );
  AOI22_X1 U558 ( .A1(data_in[3]), .A2(n1663), .B1(n829), .B2(\mem[26][3] ), 
        .ZN(n832) );
  INV_X1 U559 ( .A(n833), .ZN(n1413) );
  AOI22_X1 U560 ( .A1(data_in[4]), .A2(n1663), .B1(n829), .B2(\mem[26][4] ), 
        .ZN(n833) );
  INV_X1 U561 ( .A(n834), .ZN(n1412) );
  AOI22_X1 U562 ( .A1(data_in[5]), .A2(n1663), .B1(n829), .B2(\mem[26][5] ), 
        .ZN(n834) );
  INV_X1 U563 ( .A(n835), .ZN(n1411) );
  AOI22_X1 U564 ( .A1(data_in[6]), .A2(n1663), .B1(n829), .B2(\mem[26][6] ), 
        .ZN(n835) );
  INV_X1 U565 ( .A(n836), .ZN(n1410) );
  AOI22_X1 U566 ( .A1(data_in[7]), .A2(n1663), .B1(n829), .B2(\mem[26][7] ), 
        .ZN(n836) );
  INV_X1 U567 ( .A(n837), .ZN(n1409) );
  AOI22_X1 U568 ( .A1(data_in[0]), .A2(n1662), .B1(n838), .B2(\mem[27][0] ), 
        .ZN(n837) );
  INV_X1 U569 ( .A(n839), .ZN(n1408) );
  AOI22_X1 U570 ( .A1(data_in[1]), .A2(n1662), .B1(n838), .B2(\mem[27][1] ), 
        .ZN(n839) );
  INV_X1 U571 ( .A(n840), .ZN(n1407) );
  AOI22_X1 U572 ( .A1(data_in[2]), .A2(n1662), .B1(n838), .B2(\mem[27][2] ), 
        .ZN(n840) );
  INV_X1 U573 ( .A(n841), .ZN(n1406) );
  AOI22_X1 U574 ( .A1(data_in[3]), .A2(n1662), .B1(n838), .B2(\mem[27][3] ), 
        .ZN(n841) );
  INV_X1 U575 ( .A(n842), .ZN(n1405) );
  AOI22_X1 U576 ( .A1(data_in[4]), .A2(n1662), .B1(n838), .B2(\mem[27][4] ), 
        .ZN(n842) );
  INV_X1 U577 ( .A(n843), .ZN(n1404) );
  AOI22_X1 U578 ( .A1(data_in[5]), .A2(n1662), .B1(n838), .B2(\mem[27][5] ), 
        .ZN(n843) );
  INV_X1 U579 ( .A(n844), .ZN(n1403) );
  AOI22_X1 U580 ( .A1(data_in[6]), .A2(n1662), .B1(n838), .B2(\mem[27][6] ), 
        .ZN(n844) );
  INV_X1 U581 ( .A(n845), .ZN(n1402) );
  AOI22_X1 U582 ( .A1(data_in[7]), .A2(n1662), .B1(n838), .B2(\mem[27][7] ), 
        .ZN(n845) );
  INV_X1 U583 ( .A(n882), .ZN(n1369) );
  AOI22_X1 U584 ( .A1(data_in[0]), .A2(n1657), .B1(n883), .B2(\mem[32][0] ), 
        .ZN(n882) );
  INV_X1 U585 ( .A(n884), .ZN(n1368) );
  AOI22_X1 U586 ( .A1(data_in[1]), .A2(n1657), .B1(n883), .B2(\mem[32][1] ), 
        .ZN(n884) );
  INV_X1 U587 ( .A(n885), .ZN(n1367) );
  AOI22_X1 U588 ( .A1(data_in[2]), .A2(n1657), .B1(n883), .B2(\mem[32][2] ), 
        .ZN(n885) );
  INV_X1 U589 ( .A(n886), .ZN(n1366) );
  AOI22_X1 U590 ( .A1(data_in[3]), .A2(n1657), .B1(n883), .B2(\mem[32][3] ), 
        .ZN(n886) );
  INV_X1 U591 ( .A(n887), .ZN(n1365) );
  AOI22_X1 U592 ( .A1(data_in[4]), .A2(n1657), .B1(n883), .B2(\mem[32][4] ), 
        .ZN(n887) );
  INV_X1 U593 ( .A(n888), .ZN(n1364) );
  AOI22_X1 U594 ( .A1(data_in[5]), .A2(n1657), .B1(n883), .B2(\mem[32][5] ), 
        .ZN(n888) );
  INV_X1 U595 ( .A(n889), .ZN(n1363) );
  AOI22_X1 U596 ( .A1(data_in[6]), .A2(n1657), .B1(n883), .B2(\mem[32][6] ), 
        .ZN(n889) );
  INV_X1 U597 ( .A(n890), .ZN(n1362) );
  AOI22_X1 U598 ( .A1(data_in[7]), .A2(n1657), .B1(n883), .B2(\mem[32][7] ), 
        .ZN(n890) );
  INV_X1 U599 ( .A(n892), .ZN(n1361) );
  AOI22_X1 U600 ( .A1(data_in[0]), .A2(n1656), .B1(n893), .B2(\mem[33][0] ), 
        .ZN(n892) );
  INV_X1 U601 ( .A(n894), .ZN(n1360) );
  AOI22_X1 U602 ( .A1(data_in[1]), .A2(n1656), .B1(n893), .B2(\mem[33][1] ), 
        .ZN(n894) );
  INV_X1 U603 ( .A(n895), .ZN(n1359) );
  AOI22_X1 U604 ( .A1(data_in[2]), .A2(n1656), .B1(n893), .B2(\mem[33][2] ), 
        .ZN(n895) );
  INV_X1 U605 ( .A(n896), .ZN(n1358) );
  AOI22_X1 U606 ( .A1(data_in[3]), .A2(n1656), .B1(n893), .B2(\mem[33][3] ), 
        .ZN(n896) );
  INV_X1 U607 ( .A(n897), .ZN(n1357) );
  AOI22_X1 U608 ( .A1(data_in[4]), .A2(n1656), .B1(n893), .B2(\mem[33][4] ), 
        .ZN(n897) );
  INV_X1 U609 ( .A(n898), .ZN(n1356) );
  AOI22_X1 U610 ( .A1(data_in[5]), .A2(n1656), .B1(n893), .B2(\mem[33][5] ), 
        .ZN(n898) );
  INV_X1 U611 ( .A(n899), .ZN(n1355) );
  AOI22_X1 U612 ( .A1(data_in[6]), .A2(n1656), .B1(n893), .B2(\mem[33][6] ), 
        .ZN(n899) );
  INV_X1 U613 ( .A(n900), .ZN(n1354) );
  AOI22_X1 U614 ( .A1(data_in[7]), .A2(n1656), .B1(n893), .B2(\mem[33][7] ), 
        .ZN(n900) );
  INV_X1 U615 ( .A(n901), .ZN(n1353) );
  AOI22_X1 U616 ( .A1(data_in[0]), .A2(n1655), .B1(n902), .B2(\mem[34][0] ), 
        .ZN(n901) );
  INV_X1 U617 ( .A(n903), .ZN(n1352) );
  AOI22_X1 U618 ( .A1(data_in[1]), .A2(n1655), .B1(n902), .B2(\mem[34][1] ), 
        .ZN(n903) );
  INV_X1 U619 ( .A(n904), .ZN(n1351) );
  AOI22_X1 U620 ( .A1(data_in[2]), .A2(n1655), .B1(n902), .B2(\mem[34][2] ), 
        .ZN(n904) );
  INV_X1 U621 ( .A(n905), .ZN(n1350) );
  AOI22_X1 U622 ( .A1(data_in[3]), .A2(n1655), .B1(n902), .B2(\mem[34][3] ), 
        .ZN(n905) );
  INV_X1 U623 ( .A(n906), .ZN(n1349) );
  AOI22_X1 U624 ( .A1(data_in[4]), .A2(n1655), .B1(n902), .B2(\mem[34][4] ), 
        .ZN(n906) );
  INV_X1 U625 ( .A(n907), .ZN(n1348) );
  AOI22_X1 U626 ( .A1(data_in[5]), .A2(n1655), .B1(n902), .B2(\mem[34][5] ), 
        .ZN(n907) );
  INV_X1 U627 ( .A(n908), .ZN(n1347) );
  AOI22_X1 U628 ( .A1(data_in[6]), .A2(n1655), .B1(n902), .B2(\mem[34][6] ), 
        .ZN(n908) );
  INV_X1 U629 ( .A(n909), .ZN(n1346) );
  AOI22_X1 U630 ( .A1(data_in[7]), .A2(n1655), .B1(n902), .B2(\mem[34][7] ), 
        .ZN(n909) );
  INV_X1 U631 ( .A(n910), .ZN(n1345) );
  AOI22_X1 U632 ( .A1(data_in[0]), .A2(n1654), .B1(n911), .B2(\mem[35][0] ), 
        .ZN(n910) );
  INV_X1 U633 ( .A(n912), .ZN(n1344) );
  AOI22_X1 U634 ( .A1(data_in[1]), .A2(n1654), .B1(n911), .B2(\mem[35][1] ), 
        .ZN(n912) );
  INV_X1 U635 ( .A(n913), .ZN(n1343) );
  AOI22_X1 U636 ( .A1(data_in[2]), .A2(n1654), .B1(n911), .B2(\mem[35][2] ), 
        .ZN(n913) );
  INV_X1 U637 ( .A(n914), .ZN(n1342) );
  AOI22_X1 U638 ( .A1(data_in[3]), .A2(n1654), .B1(n911), .B2(\mem[35][3] ), 
        .ZN(n914) );
  INV_X1 U639 ( .A(n915), .ZN(n1341) );
  AOI22_X1 U640 ( .A1(data_in[4]), .A2(n1654), .B1(n911), .B2(\mem[35][4] ), 
        .ZN(n915) );
  INV_X1 U641 ( .A(n916), .ZN(n1340) );
  AOI22_X1 U642 ( .A1(data_in[5]), .A2(n1654), .B1(n911), .B2(\mem[35][5] ), 
        .ZN(n916) );
  INV_X1 U643 ( .A(n917), .ZN(n1339) );
  AOI22_X1 U644 ( .A1(data_in[6]), .A2(n1654), .B1(n911), .B2(\mem[35][6] ), 
        .ZN(n917) );
  INV_X1 U645 ( .A(n918), .ZN(n1338) );
  AOI22_X1 U646 ( .A1(data_in[7]), .A2(n1654), .B1(n911), .B2(\mem[35][7] ), 
        .ZN(n918) );
  INV_X1 U647 ( .A(n955), .ZN(n1305) );
  AOI22_X1 U648 ( .A1(data_in[0]), .A2(n1649), .B1(n956), .B2(\mem[40][0] ), 
        .ZN(n955) );
  INV_X1 U649 ( .A(n957), .ZN(n1304) );
  AOI22_X1 U650 ( .A1(data_in[1]), .A2(n1649), .B1(n956), .B2(\mem[40][1] ), 
        .ZN(n957) );
  INV_X1 U651 ( .A(n958), .ZN(n1303) );
  AOI22_X1 U652 ( .A1(data_in[2]), .A2(n1649), .B1(n956), .B2(\mem[40][2] ), 
        .ZN(n958) );
  INV_X1 U653 ( .A(n959), .ZN(n1302) );
  AOI22_X1 U654 ( .A1(data_in[3]), .A2(n1649), .B1(n956), .B2(\mem[40][3] ), 
        .ZN(n959) );
  INV_X1 U655 ( .A(n960), .ZN(n1301) );
  AOI22_X1 U656 ( .A1(data_in[4]), .A2(n1649), .B1(n956), .B2(\mem[40][4] ), 
        .ZN(n960) );
  INV_X1 U657 ( .A(n961), .ZN(n1300) );
  AOI22_X1 U658 ( .A1(data_in[5]), .A2(n1649), .B1(n956), .B2(\mem[40][5] ), 
        .ZN(n961) );
  INV_X1 U659 ( .A(n962), .ZN(n1299) );
  AOI22_X1 U660 ( .A1(data_in[6]), .A2(n1649), .B1(n956), .B2(\mem[40][6] ), 
        .ZN(n962) );
  INV_X1 U661 ( .A(n963), .ZN(n1298) );
  AOI22_X1 U662 ( .A1(data_in[7]), .A2(n1649), .B1(n956), .B2(\mem[40][7] ), 
        .ZN(n963) );
  INV_X1 U663 ( .A(n965), .ZN(n1297) );
  AOI22_X1 U664 ( .A1(data_in[0]), .A2(n1648), .B1(n966), .B2(\mem[41][0] ), 
        .ZN(n965) );
  INV_X1 U665 ( .A(n967), .ZN(n1296) );
  AOI22_X1 U666 ( .A1(data_in[1]), .A2(n1648), .B1(n966), .B2(\mem[41][1] ), 
        .ZN(n967) );
  INV_X1 U667 ( .A(n968), .ZN(n1295) );
  AOI22_X1 U668 ( .A1(data_in[2]), .A2(n1648), .B1(n966), .B2(\mem[41][2] ), 
        .ZN(n968) );
  INV_X1 U669 ( .A(n969), .ZN(n1294) );
  AOI22_X1 U670 ( .A1(data_in[3]), .A2(n1648), .B1(n966), .B2(\mem[41][3] ), 
        .ZN(n969) );
  INV_X1 U671 ( .A(n970), .ZN(n1293) );
  AOI22_X1 U672 ( .A1(data_in[4]), .A2(n1648), .B1(n966), .B2(\mem[41][4] ), 
        .ZN(n970) );
  INV_X1 U673 ( .A(n971), .ZN(n1292) );
  AOI22_X1 U674 ( .A1(data_in[5]), .A2(n1648), .B1(n966), .B2(\mem[41][5] ), 
        .ZN(n971) );
  INV_X1 U675 ( .A(n972), .ZN(n1291) );
  AOI22_X1 U676 ( .A1(data_in[6]), .A2(n1648), .B1(n966), .B2(\mem[41][6] ), 
        .ZN(n972) );
  INV_X1 U677 ( .A(n973), .ZN(n1290) );
  AOI22_X1 U678 ( .A1(data_in[7]), .A2(n1648), .B1(n966), .B2(\mem[41][7] ), 
        .ZN(n973) );
  INV_X1 U679 ( .A(n974), .ZN(n1289) );
  AOI22_X1 U680 ( .A1(data_in[0]), .A2(n1647), .B1(n975), .B2(\mem[42][0] ), 
        .ZN(n974) );
  INV_X1 U681 ( .A(n976), .ZN(n1288) );
  AOI22_X1 U682 ( .A1(data_in[1]), .A2(n1647), .B1(n975), .B2(\mem[42][1] ), 
        .ZN(n976) );
  INV_X1 U683 ( .A(n977), .ZN(n1287) );
  AOI22_X1 U684 ( .A1(data_in[2]), .A2(n1647), .B1(n975), .B2(\mem[42][2] ), 
        .ZN(n977) );
  INV_X1 U685 ( .A(n978), .ZN(n1286) );
  AOI22_X1 U686 ( .A1(data_in[3]), .A2(n1647), .B1(n975), .B2(\mem[42][3] ), 
        .ZN(n978) );
  INV_X1 U687 ( .A(n979), .ZN(n1285) );
  AOI22_X1 U688 ( .A1(data_in[4]), .A2(n1647), .B1(n975), .B2(\mem[42][4] ), 
        .ZN(n979) );
  INV_X1 U689 ( .A(n980), .ZN(n1284) );
  AOI22_X1 U690 ( .A1(data_in[5]), .A2(n1647), .B1(n975), .B2(\mem[42][5] ), 
        .ZN(n980) );
  INV_X1 U691 ( .A(n981), .ZN(n1283) );
  AOI22_X1 U692 ( .A1(data_in[6]), .A2(n1647), .B1(n975), .B2(\mem[42][6] ), 
        .ZN(n981) );
  INV_X1 U693 ( .A(n982), .ZN(n1282) );
  AOI22_X1 U694 ( .A1(data_in[7]), .A2(n1647), .B1(n975), .B2(\mem[42][7] ), 
        .ZN(n982) );
  INV_X1 U695 ( .A(n983), .ZN(n1281) );
  AOI22_X1 U696 ( .A1(data_in[0]), .A2(n1646), .B1(n984), .B2(\mem[43][0] ), 
        .ZN(n983) );
  INV_X1 U697 ( .A(n985), .ZN(n1280) );
  AOI22_X1 U698 ( .A1(data_in[1]), .A2(n1646), .B1(n984), .B2(\mem[43][1] ), 
        .ZN(n985) );
  INV_X1 U699 ( .A(n986), .ZN(n1279) );
  AOI22_X1 U700 ( .A1(data_in[2]), .A2(n1646), .B1(n984), .B2(\mem[43][2] ), 
        .ZN(n986) );
  INV_X1 U701 ( .A(n987), .ZN(n1278) );
  AOI22_X1 U702 ( .A1(data_in[3]), .A2(n1646), .B1(n984), .B2(\mem[43][3] ), 
        .ZN(n987) );
  INV_X1 U703 ( .A(n988), .ZN(n1277) );
  AOI22_X1 U704 ( .A1(data_in[4]), .A2(n1646), .B1(n984), .B2(\mem[43][4] ), 
        .ZN(n988) );
  INV_X1 U705 ( .A(n989), .ZN(n1276) );
  AOI22_X1 U706 ( .A1(data_in[5]), .A2(n1646), .B1(n984), .B2(\mem[43][5] ), 
        .ZN(n989) );
  INV_X1 U707 ( .A(n990), .ZN(n1275) );
  AOI22_X1 U708 ( .A1(data_in[6]), .A2(n1646), .B1(n984), .B2(\mem[43][6] ), 
        .ZN(n990) );
  INV_X1 U709 ( .A(n991), .ZN(n1274) );
  AOI22_X1 U710 ( .A1(data_in[7]), .A2(n1646), .B1(n984), .B2(\mem[43][7] ), 
        .ZN(n991) );
  INV_X1 U711 ( .A(n1028), .ZN(n1241) );
  AOI22_X1 U712 ( .A1(data_in[0]), .A2(n1641), .B1(n1029), .B2(\mem[48][0] ), 
        .ZN(n1028) );
  INV_X1 U713 ( .A(n1030), .ZN(n1240) );
  AOI22_X1 U714 ( .A1(data_in[1]), .A2(n1641), .B1(n1029), .B2(\mem[48][1] ), 
        .ZN(n1030) );
  INV_X1 U715 ( .A(n1031), .ZN(n1239) );
  AOI22_X1 U716 ( .A1(data_in[2]), .A2(n1641), .B1(n1029), .B2(\mem[48][2] ), 
        .ZN(n1031) );
  INV_X1 U717 ( .A(n1032), .ZN(n1238) );
  AOI22_X1 U718 ( .A1(data_in[3]), .A2(n1641), .B1(n1029), .B2(\mem[48][3] ), 
        .ZN(n1032) );
  INV_X1 U719 ( .A(n1033), .ZN(n1237) );
  AOI22_X1 U720 ( .A1(data_in[4]), .A2(n1641), .B1(n1029), .B2(\mem[48][4] ), 
        .ZN(n1033) );
  INV_X1 U721 ( .A(n1034), .ZN(n1236) );
  AOI22_X1 U722 ( .A1(data_in[5]), .A2(n1641), .B1(n1029), .B2(\mem[48][5] ), 
        .ZN(n1034) );
  INV_X1 U723 ( .A(n1035), .ZN(n1235) );
  AOI22_X1 U724 ( .A1(data_in[6]), .A2(n1641), .B1(n1029), .B2(\mem[48][6] ), 
        .ZN(n1035) );
  INV_X1 U725 ( .A(n1036), .ZN(n1234) );
  AOI22_X1 U726 ( .A1(data_in[7]), .A2(n1641), .B1(n1029), .B2(\mem[48][7] ), 
        .ZN(n1036) );
  INV_X1 U727 ( .A(n1038), .ZN(n1233) );
  AOI22_X1 U728 ( .A1(data_in[0]), .A2(n1640), .B1(n1039), .B2(\mem[49][0] ), 
        .ZN(n1038) );
  INV_X1 U729 ( .A(n1040), .ZN(n1232) );
  AOI22_X1 U730 ( .A1(data_in[1]), .A2(n1640), .B1(n1039), .B2(\mem[49][1] ), 
        .ZN(n1040) );
  INV_X1 U731 ( .A(n1041), .ZN(n1231) );
  AOI22_X1 U732 ( .A1(data_in[2]), .A2(n1640), .B1(n1039), .B2(\mem[49][2] ), 
        .ZN(n1041) );
  INV_X1 U733 ( .A(n1042), .ZN(n1230) );
  AOI22_X1 U734 ( .A1(data_in[3]), .A2(n1640), .B1(n1039), .B2(\mem[49][3] ), 
        .ZN(n1042) );
  INV_X1 U735 ( .A(n1043), .ZN(n1229) );
  AOI22_X1 U736 ( .A1(data_in[4]), .A2(n1640), .B1(n1039), .B2(\mem[49][4] ), 
        .ZN(n1043) );
  INV_X1 U737 ( .A(n1044), .ZN(n1228) );
  AOI22_X1 U738 ( .A1(data_in[5]), .A2(n1640), .B1(n1039), .B2(\mem[49][5] ), 
        .ZN(n1044) );
  INV_X1 U739 ( .A(n1045), .ZN(n1227) );
  AOI22_X1 U740 ( .A1(data_in[6]), .A2(n1640), .B1(n1039), .B2(\mem[49][6] ), 
        .ZN(n1045) );
  INV_X1 U741 ( .A(n1046), .ZN(n1226) );
  AOI22_X1 U742 ( .A1(data_in[7]), .A2(n1640), .B1(n1039), .B2(\mem[49][7] ), 
        .ZN(n1046) );
  INV_X1 U743 ( .A(n1047), .ZN(n1225) );
  AOI22_X1 U744 ( .A1(data_in[0]), .A2(n1639), .B1(n1048), .B2(\mem[50][0] ), 
        .ZN(n1047) );
  INV_X1 U745 ( .A(n1049), .ZN(n1224) );
  AOI22_X1 U746 ( .A1(data_in[1]), .A2(n1639), .B1(n1048), .B2(\mem[50][1] ), 
        .ZN(n1049) );
  INV_X1 U747 ( .A(n1050), .ZN(n1223) );
  AOI22_X1 U748 ( .A1(data_in[2]), .A2(n1639), .B1(n1048), .B2(\mem[50][2] ), 
        .ZN(n1050) );
  INV_X1 U749 ( .A(n1051), .ZN(n1222) );
  AOI22_X1 U750 ( .A1(data_in[3]), .A2(n1639), .B1(n1048), .B2(\mem[50][3] ), 
        .ZN(n1051) );
  INV_X1 U751 ( .A(n1052), .ZN(n1221) );
  AOI22_X1 U752 ( .A1(data_in[4]), .A2(n1639), .B1(n1048), .B2(\mem[50][4] ), 
        .ZN(n1052) );
  INV_X1 U753 ( .A(n1053), .ZN(n1220) );
  AOI22_X1 U754 ( .A1(data_in[5]), .A2(n1639), .B1(n1048), .B2(\mem[50][5] ), 
        .ZN(n1053) );
  INV_X1 U755 ( .A(n1054), .ZN(n1219) );
  AOI22_X1 U756 ( .A1(data_in[6]), .A2(n1639), .B1(n1048), .B2(\mem[50][6] ), 
        .ZN(n1054) );
  INV_X1 U757 ( .A(n1055), .ZN(n1218) );
  AOI22_X1 U758 ( .A1(data_in[7]), .A2(n1639), .B1(n1048), .B2(\mem[50][7] ), 
        .ZN(n1055) );
  INV_X1 U759 ( .A(n1056), .ZN(n1217) );
  AOI22_X1 U760 ( .A1(data_in[0]), .A2(n1638), .B1(n1057), .B2(\mem[51][0] ), 
        .ZN(n1056) );
  INV_X1 U761 ( .A(n1058), .ZN(n1216) );
  AOI22_X1 U762 ( .A1(data_in[1]), .A2(n1638), .B1(n1057), .B2(\mem[51][1] ), 
        .ZN(n1058) );
  INV_X1 U763 ( .A(n1059), .ZN(n1215) );
  AOI22_X1 U764 ( .A1(data_in[2]), .A2(n1638), .B1(n1057), .B2(\mem[51][2] ), 
        .ZN(n1059) );
  INV_X1 U765 ( .A(n1060), .ZN(n1214) );
  AOI22_X1 U766 ( .A1(data_in[3]), .A2(n1638), .B1(n1057), .B2(\mem[51][3] ), 
        .ZN(n1060) );
  INV_X1 U767 ( .A(n1061), .ZN(n1213) );
  AOI22_X1 U768 ( .A1(data_in[4]), .A2(n1638), .B1(n1057), .B2(\mem[51][4] ), 
        .ZN(n1061) );
  INV_X1 U769 ( .A(n1062), .ZN(n1212) );
  AOI22_X1 U770 ( .A1(data_in[5]), .A2(n1638), .B1(n1057), .B2(\mem[51][5] ), 
        .ZN(n1062) );
  INV_X1 U771 ( .A(n1063), .ZN(n1211) );
  AOI22_X1 U772 ( .A1(data_in[6]), .A2(n1638), .B1(n1057), .B2(\mem[51][6] ), 
        .ZN(n1063) );
  INV_X1 U773 ( .A(n1064), .ZN(n1210) );
  AOI22_X1 U774 ( .A1(data_in[7]), .A2(n1638), .B1(n1057), .B2(\mem[51][7] ), 
        .ZN(n1064) );
  INV_X1 U775 ( .A(n1101), .ZN(n1177) );
  AOI22_X1 U776 ( .A1(data_in[0]), .A2(n1633), .B1(n1102), .B2(\mem[56][0] ), 
        .ZN(n1101) );
  INV_X1 U777 ( .A(n1103), .ZN(n1176) );
  AOI22_X1 U778 ( .A1(data_in[1]), .A2(n1633), .B1(n1102), .B2(\mem[56][1] ), 
        .ZN(n1103) );
  INV_X1 U779 ( .A(n1104), .ZN(n1175) );
  AOI22_X1 U780 ( .A1(data_in[2]), .A2(n1633), .B1(n1102), .B2(\mem[56][2] ), 
        .ZN(n1104) );
  INV_X1 U781 ( .A(n1105), .ZN(n1174) );
  AOI22_X1 U782 ( .A1(data_in[3]), .A2(n1633), .B1(n1102), .B2(\mem[56][3] ), 
        .ZN(n1105) );
  INV_X1 U783 ( .A(n1106), .ZN(n581) );
  AOI22_X1 U784 ( .A1(data_in[4]), .A2(n1633), .B1(n1102), .B2(\mem[56][4] ), 
        .ZN(n1106) );
  INV_X1 U785 ( .A(n1107), .ZN(n580) );
  AOI22_X1 U786 ( .A1(data_in[5]), .A2(n1633), .B1(n1102), .B2(\mem[56][5] ), 
        .ZN(n1107) );
  INV_X1 U787 ( .A(n1108), .ZN(n579) );
  AOI22_X1 U788 ( .A1(data_in[6]), .A2(n1633), .B1(n1102), .B2(\mem[56][6] ), 
        .ZN(n1108) );
  INV_X1 U789 ( .A(n1109), .ZN(n578) );
  AOI22_X1 U790 ( .A1(data_in[7]), .A2(n1633), .B1(n1102), .B2(\mem[56][7] ), 
        .ZN(n1109) );
  INV_X1 U791 ( .A(n1111), .ZN(n577) );
  AOI22_X1 U792 ( .A1(data_in[0]), .A2(n1632), .B1(n1112), .B2(\mem[57][0] ), 
        .ZN(n1111) );
  INV_X1 U793 ( .A(n1113), .ZN(n576) );
  AOI22_X1 U794 ( .A1(data_in[1]), .A2(n1632), .B1(n1112), .B2(\mem[57][1] ), 
        .ZN(n1113) );
  INV_X1 U795 ( .A(n1114), .ZN(n575) );
  AOI22_X1 U796 ( .A1(data_in[2]), .A2(n1632), .B1(n1112), .B2(\mem[57][2] ), 
        .ZN(n1114) );
  INV_X1 U797 ( .A(n1115), .ZN(n574) );
  AOI22_X1 U798 ( .A1(data_in[3]), .A2(n1632), .B1(n1112), .B2(\mem[57][3] ), 
        .ZN(n1115) );
  INV_X1 U799 ( .A(n1116), .ZN(n573) );
  AOI22_X1 U800 ( .A1(data_in[4]), .A2(n1632), .B1(n1112), .B2(\mem[57][4] ), 
        .ZN(n1116) );
  INV_X1 U801 ( .A(n1117), .ZN(n572) );
  AOI22_X1 U802 ( .A1(data_in[5]), .A2(n1632), .B1(n1112), .B2(\mem[57][5] ), 
        .ZN(n1117) );
  INV_X1 U803 ( .A(n1118), .ZN(n571) );
  AOI22_X1 U804 ( .A1(data_in[6]), .A2(n1632), .B1(n1112), .B2(\mem[57][6] ), 
        .ZN(n1118) );
  INV_X1 U805 ( .A(n1119), .ZN(n570) );
  AOI22_X1 U806 ( .A1(data_in[7]), .A2(n1632), .B1(n1112), .B2(\mem[57][7] ), 
        .ZN(n1119) );
  INV_X1 U807 ( .A(n1120), .ZN(n569) );
  AOI22_X1 U808 ( .A1(data_in[0]), .A2(n1631), .B1(n1121), .B2(\mem[58][0] ), 
        .ZN(n1120) );
  INV_X1 U809 ( .A(n1122), .ZN(n568) );
  AOI22_X1 U810 ( .A1(data_in[1]), .A2(n1631), .B1(n1121), .B2(\mem[58][1] ), 
        .ZN(n1122) );
  INV_X1 U811 ( .A(n1123), .ZN(n567) );
  AOI22_X1 U812 ( .A1(data_in[2]), .A2(n1631), .B1(n1121), .B2(\mem[58][2] ), 
        .ZN(n1123) );
  INV_X1 U813 ( .A(n1124), .ZN(n566) );
  AOI22_X1 U814 ( .A1(data_in[3]), .A2(n1631), .B1(n1121), .B2(\mem[58][3] ), 
        .ZN(n1124) );
  INV_X1 U815 ( .A(n1125), .ZN(n565) );
  AOI22_X1 U816 ( .A1(data_in[4]), .A2(n1631), .B1(n1121), .B2(\mem[58][4] ), 
        .ZN(n1125) );
  INV_X1 U817 ( .A(n1126), .ZN(n564) );
  AOI22_X1 U818 ( .A1(data_in[5]), .A2(n1631), .B1(n1121), .B2(\mem[58][5] ), 
        .ZN(n1126) );
  INV_X1 U819 ( .A(n1127), .ZN(n563) );
  AOI22_X1 U820 ( .A1(data_in[6]), .A2(n1631), .B1(n1121), .B2(\mem[58][6] ), 
        .ZN(n1127) );
  INV_X1 U821 ( .A(n1128), .ZN(n562) );
  AOI22_X1 U822 ( .A1(data_in[7]), .A2(n1631), .B1(n1121), .B2(\mem[58][7] ), 
        .ZN(n1128) );
  INV_X1 U823 ( .A(n1129), .ZN(n561) );
  AOI22_X1 U824 ( .A1(data_in[0]), .A2(n1630), .B1(n1130), .B2(\mem[59][0] ), 
        .ZN(n1129) );
  INV_X1 U825 ( .A(n1131), .ZN(n560) );
  AOI22_X1 U826 ( .A1(data_in[1]), .A2(n1630), .B1(n1130), .B2(\mem[59][1] ), 
        .ZN(n1131) );
  INV_X1 U827 ( .A(n1132), .ZN(n559) );
  AOI22_X1 U828 ( .A1(data_in[2]), .A2(n1630), .B1(n1130), .B2(\mem[59][2] ), 
        .ZN(n1132) );
  INV_X1 U829 ( .A(n1133), .ZN(n558) );
  AOI22_X1 U830 ( .A1(data_in[3]), .A2(n1630), .B1(n1130), .B2(\mem[59][3] ), 
        .ZN(n1133) );
  INV_X1 U831 ( .A(n1134), .ZN(n557) );
  AOI22_X1 U832 ( .A1(data_in[4]), .A2(n1630), .B1(n1130), .B2(\mem[59][4] ), 
        .ZN(n1134) );
  INV_X1 U833 ( .A(n1135), .ZN(n556) );
  AOI22_X1 U834 ( .A1(data_in[5]), .A2(n1630), .B1(n1130), .B2(\mem[59][5] ), 
        .ZN(n1135) );
  INV_X1 U835 ( .A(n1136), .ZN(n555) );
  AOI22_X1 U836 ( .A1(data_in[6]), .A2(n1630), .B1(n1130), .B2(\mem[59][6] ), 
        .ZN(n1136) );
  INV_X1 U837 ( .A(n1137), .ZN(n554) );
  AOI22_X1 U838 ( .A1(data_in[7]), .A2(n1630), .B1(n1130), .B2(\mem[59][7] ), 
        .ZN(n1137) );
  INV_X1 U839 ( .A(n709), .ZN(n1521) );
  AOI22_X1 U840 ( .A1(data_in[0]), .A2(n1676), .B1(n710), .B2(\mem[13][0] ), 
        .ZN(n709) );
  INV_X1 U841 ( .A(n711), .ZN(n1520) );
  AOI22_X1 U842 ( .A1(data_in[1]), .A2(n1676), .B1(n710), .B2(\mem[13][1] ), 
        .ZN(n711) );
  INV_X1 U843 ( .A(n712), .ZN(n1519) );
  AOI22_X1 U844 ( .A1(data_in[2]), .A2(n1676), .B1(n710), .B2(\mem[13][2] ), 
        .ZN(n712) );
  INV_X1 U845 ( .A(n713), .ZN(n1518) );
  AOI22_X1 U846 ( .A1(data_in[3]), .A2(n1676), .B1(n710), .B2(\mem[13][3] ), 
        .ZN(n713) );
  INV_X1 U847 ( .A(n714), .ZN(n1517) );
  AOI22_X1 U848 ( .A1(data_in[4]), .A2(n1676), .B1(n710), .B2(\mem[13][4] ), 
        .ZN(n714) );
  INV_X1 U849 ( .A(n715), .ZN(n1516) );
  AOI22_X1 U850 ( .A1(data_in[5]), .A2(n1676), .B1(n710), .B2(\mem[13][5] ), 
        .ZN(n715) );
  INV_X1 U851 ( .A(n716), .ZN(n1515) );
  AOI22_X1 U852 ( .A1(data_in[6]), .A2(n1676), .B1(n710), .B2(\mem[13][6] ), 
        .ZN(n716) );
  INV_X1 U853 ( .A(n717), .ZN(n1514) );
  AOI22_X1 U854 ( .A1(data_in[7]), .A2(n1676), .B1(n710), .B2(\mem[13][7] ), 
        .ZN(n717) );
  INV_X1 U855 ( .A(n727), .ZN(n1505) );
  AOI22_X1 U856 ( .A1(data_in[0]), .A2(n1674), .B1(n728), .B2(\mem[15][0] ), 
        .ZN(n727) );
  INV_X1 U857 ( .A(n729), .ZN(n1504) );
  AOI22_X1 U858 ( .A1(data_in[1]), .A2(n1674), .B1(n728), .B2(\mem[15][1] ), 
        .ZN(n729) );
  INV_X1 U859 ( .A(n730), .ZN(n1503) );
  AOI22_X1 U860 ( .A1(data_in[2]), .A2(n1674), .B1(n728), .B2(\mem[15][2] ), 
        .ZN(n730) );
  INV_X1 U861 ( .A(n731), .ZN(n1502) );
  AOI22_X1 U862 ( .A1(data_in[3]), .A2(n1674), .B1(n728), .B2(\mem[15][3] ), 
        .ZN(n731) );
  INV_X1 U863 ( .A(n732), .ZN(n1501) );
  AOI22_X1 U864 ( .A1(data_in[4]), .A2(n1674), .B1(n728), .B2(\mem[15][4] ), 
        .ZN(n732) );
  INV_X1 U865 ( .A(n733), .ZN(n1500) );
  AOI22_X1 U866 ( .A1(data_in[5]), .A2(n1674), .B1(n728), .B2(\mem[15][5] ), 
        .ZN(n733) );
  INV_X1 U867 ( .A(n734), .ZN(n1499) );
  AOI22_X1 U868 ( .A1(data_in[6]), .A2(n1674), .B1(n728), .B2(\mem[15][6] ), 
        .ZN(n734) );
  INV_X1 U869 ( .A(n735), .ZN(n1498) );
  AOI22_X1 U870 ( .A1(data_in[7]), .A2(n1674), .B1(n728), .B2(\mem[15][7] ), 
        .ZN(n735) );
  INV_X1 U871 ( .A(n782), .ZN(n1457) );
  AOI22_X1 U872 ( .A1(data_in[0]), .A2(n1668), .B1(n783), .B2(\mem[21][0] ), 
        .ZN(n782) );
  INV_X1 U873 ( .A(n784), .ZN(n1456) );
  AOI22_X1 U874 ( .A1(data_in[1]), .A2(n1668), .B1(n783), .B2(\mem[21][1] ), 
        .ZN(n784) );
  INV_X1 U875 ( .A(n785), .ZN(n1455) );
  AOI22_X1 U876 ( .A1(data_in[2]), .A2(n1668), .B1(n783), .B2(\mem[21][2] ), 
        .ZN(n785) );
  INV_X1 U877 ( .A(n786), .ZN(n1454) );
  AOI22_X1 U878 ( .A1(data_in[3]), .A2(n1668), .B1(n783), .B2(\mem[21][3] ), 
        .ZN(n786) );
  INV_X1 U879 ( .A(n787), .ZN(n1453) );
  AOI22_X1 U880 ( .A1(data_in[4]), .A2(n1668), .B1(n783), .B2(\mem[21][4] ), 
        .ZN(n787) );
  INV_X1 U881 ( .A(n788), .ZN(n1452) );
  AOI22_X1 U882 ( .A1(data_in[5]), .A2(n1668), .B1(n783), .B2(\mem[21][5] ), 
        .ZN(n788) );
  INV_X1 U883 ( .A(n789), .ZN(n1451) );
  AOI22_X1 U884 ( .A1(data_in[6]), .A2(n1668), .B1(n783), .B2(\mem[21][6] ), 
        .ZN(n789) );
  INV_X1 U885 ( .A(n790), .ZN(n1450) );
  AOI22_X1 U886 ( .A1(data_in[7]), .A2(n1668), .B1(n783), .B2(\mem[21][7] ), 
        .ZN(n790) );
  INV_X1 U887 ( .A(n800), .ZN(n1441) );
  AOI22_X1 U888 ( .A1(data_in[0]), .A2(n1666), .B1(n801), .B2(\mem[23][0] ), 
        .ZN(n800) );
  INV_X1 U889 ( .A(n802), .ZN(n1440) );
  AOI22_X1 U890 ( .A1(data_in[1]), .A2(n1666), .B1(n801), .B2(\mem[23][1] ), 
        .ZN(n802) );
  INV_X1 U891 ( .A(n803), .ZN(n1439) );
  AOI22_X1 U892 ( .A1(data_in[2]), .A2(n1666), .B1(n801), .B2(\mem[23][2] ), 
        .ZN(n803) );
  INV_X1 U893 ( .A(n804), .ZN(n1438) );
  AOI22_X1 U894 ( .A1(data_in[3]), .A2(n1666), .B1(n801), .B2(\mem[23][3] ), 
        .ZN(n804) );
  INV_X1 U895 ( .A(n805), .ZN(n1437) );
  AOI22_X1 U896 ( .A1(data_in[4]), .A2(n1666), .B1(n801), .B2(\mem[23][4] ), 
        .ZN(n805) );
  INV_X1 U897 ( .A(n806), .ZN(n1436) );
  AOI22_X1 U898 ( .A1(data_in[5]), .A2(n1666), .B1(n801), .B2(\mem[23][5] ), 
        .ZN(n806) );
  INV_X1 U899 ( .A(n807), .ZN(n1435) );
  AOI22_X1 U900 ( .A1(data_in[6]), .A2(n1666), .B1(n801), .B2(\mem[23][6] ), 
        .ZN(n807) );
  INV_X1 U901 ( .A(n808), .ZN(n1434) );
  AOI22_X1 U902 ( .A1(data_in[7]), .A2(n1666), .B1(n801), .B2(\mem[23][7] ), 
        .ZN(n808) );
  INV_X1 U903 ( .A(n855), .ZN(n1393) );
  AOI22_X1 U904 ( .A1(data_in[0]), .A2(n1660), .B1(n856), .B2(\mem[29][0] ), 
        .ZN(n855) );
  INV_X1 U905 ( .A(n857), .ZN(n1392) );
  AOI22_X1 U906 ( .A1(data_in[1]), .A2(n1660), .B1(n856), .B2(\mem[29][1] ), 
        .ZN(n857) );
  INV_X1 U907 ( .A(n858), .ZN(n1391) );
  AOI22_X1 U908 ( .A1(data_in[2]), .A2(n1660), .B1(n856), .B2(\mem[29][2] ), 
        .ZN(n858) );
  INV_X1 U909 ( .A(n859), .ZN(n1390) );
  AOI22_X1 U910 ( .A1(data_in[3]), .A2(n1660), .B1(n856), .B2(\mem[29][3] ), 
        .ZN(n859) );
  INV_X1 U911 ( .A(n860), .ZN(n1389) );
  AOI22_X1 U912 ( .A1(data_in[4]), .A2(n1660), .B1(n856), .B2(\mem[29][4] ), 
        .ZN(n860) );
  INV_X1 U913 ( .A(n861), .ZN(n1388) );
  AOI22_X1 U914 ( .A1(data_in[5]), .A2(n1660), .B1(n856), .B2(\mem[29][5] ), 
        .ZN(n861) );
  INV_X1 U915 ( .A(n862), .ZN(n1387) );
  AOI22_X1 U916 ( .A1(data_in[6]), .A2(n1660), .B1(n856), .B2(\mem[29][6] ), 
        .ZN(n862) );
  INV_X1 U917 ( .A(n863), .ZN(n1386) );
  AOI22_X1 U918 ( .A1(data_in[7]), .A2(n1660), .B1(n856), .B2(\mem[29][7] ), 
        .ZN(n863) );
  INV_X1 U919 ( .A(n873), .ZN(n1377) );
  AOI22_X1 U920 ( .A1(data_in[0]), .A2(n1658), .B1(n874), .B2(\mem[31][0] ), 
        .ZN(n873) );
  INV_X1 U921 ( .A(n875), .ZN(n1376) );
  AOI22_X1 U922 ( .A1(data_in[1]), .A2(n1658), .B1(n874), .B2(\mem[31][1] ), 
        .ZN(n875) );
  INV_X1 U923 ( .A(n876), .ZN(n1375) );
  AOI22_X1 U924 ( .A1(data_in[2]), .A2(n1658), .B1(n874), .B2(\mem[31][2] ), 
        .ZN(n876) );
  INV_X1 U925 ( .A(n877), .ZN(n1374) );
  AOI22_X1 U926 ( .A1(data_in[3]), .A2(n1658), .B1(n874), .B2(\mem[31][3] ), 
        .ZN(n877) );
  INV_X1 U927 ( .A(n878), .ZN(n1373) );
  AOI22_X1 U928 ( .A1(data_in[4]), .A2(n1658), .B1(n874), .B2(\mem[31][4] ), 
        .ZN(n878) );
  INV_X1 U929 ( .A(n879), .ZN(n1372) );
  AOI22_X1 U930 ( .A1(data_in[5]), .A2(n1658), .B1(n874), .B2(\mem[31][5] ), 
        .ZN(n879) );
  INV_X1 U931 ( .A(n880), .ZN(n1371) );
  AOI22_X1 U932 ( .A1(data_in[6]), .A2(n1658), .B1(n874), .B2(\mem[31][6] ), 
        .ZN(n880) );
  INV_X1 U933 ( .A(n881), .ZN(n1370) );
  AOI22_X1 U934 ( .A1(data_in[7]), .A2(n1658), .B1(n874), .B2(\mem[31][7] ), 
        .ZN(n881) );
  INV_X1 U935 ( .A(n928), .ZN(n1329) );
  AOI22_X1 U936 ( .A1(data_in[0]), .A2(n1652), .B1(n929), .B2(\mem[37][0] ), 
        .ZN(n928) );
  INV_X1 U937 ( .A(n930), .ZN(n1328) );
  AOI22_X1 U938 ( .A1(data_in[1]), .A2(n1652), .B1(n929), .B2(\mem[37][1] ), 
        .ZN(n930) );
  INV_X1 U939 ( .A(n931), .ZN(n1327) );
  AOI22_X1 U940 ( .A1(data_in[2]), .A2(n1652), .B1(n929), .B2(\mem[37][2] ), 
        .ZN(n931) );
  INV_X1 U941 ( .A(n932), .ZN(n1326) );
  AOI22_X1 U942 ( .A1(data_in[3]), .A2(n1652), .B1(n929), .B2(\mem[37][3] ), 
        .ZN(n932) );
  INV_X1 U943 ( .A(n933), .ZN(n1325) );
  AOI22_X1 U944 ( .A1(data_in[4]), .A2(n1652), .B1(n929), .B2(\mem[37][4] ), 
        .ZN(n933) );
  INV_X1 U945 ( .A(n934), .ZN(n1324) );
  AOI22_X1 U946 ( .A1(data_in[5]), .A2(n1652), .B1(n929), .B2(\mem[37][5] ), 
        .ZN(n934) );
  INV_X1 U947 ( .A(n935), .ZN(n1323) );
  AOI22_X1 U948 ( .A1(data_in[6]), .A2(n1652), .B1(n929), .B2(\mem[37][6] ), 
        .ZN(n935) );
  INV_X1 U949 ( .A(n936), .ZN(n1322) );
  AOI22_X1 U950 ( .A1(data_in[7]), .A2(n1652), .B1(n929), .B2(\mem[37][7] ), 
        .ZN(n936) );
  INV_X1 U951 ( .A(n946), .ZN(n1313) );
  AOI22_X1 U952 ( .A1(data_in[0]), .A2(n1650), .B1(n947), .B2(\mem[39][0] ), 
        .ZN(n946) );
  INV_X1 U953 ( .A(n948), .ZN(n1312) );
  AOI22_X1 U954 ( .A1(data_in[1]), .A2(n1650), .B1(n947), .B2(\mem[39][1] ), 
        .ZN(n948) );
  INV_X1 U955 ( .A(n949), .ZN(n1311) );
  AOI22_X1 U956 ( .A1(data_in[2]), .A2(n1650), .B1(n947), .B2(\mem[39][2] ), 
        .ZN(n949) );
  INV_X1 U957 ( .A(n950), .ZN(n1310) );
  AOI22_X1 U958 ( .A1(data_in[3]), .A2(n1650), .B1(n947), .B2(\mem[39][3] ), 
        .ZN(n950) );
  INV_X1 U959 ( .A(n951), .ZN(n1309) );
  AOI22_X1 U960 ( .A1(data_in[4]), .A2(n1650), .B1(n947), .B2(\mem[39][4] ), 
        .ZN(n951) );
  INV_X1 U961 ( .A(n952), .ZN(n1308) );
  AOI22_X1 U962 ( .A1(data_in[5]), .A2(n1650), .B1(n947), .B2(\mem[39][5] ), 
        .ZN(n952) );
  INV_X1 U963 ( .A(n953), .ZN(n1307) );
  AOI22_X1 U964 ( .A1(data_in[6]), .A2(n1650), .B1(n947), .B2(\mem[39][6] ), 
        .ZN(n953) );
  INV_X1 U965 ( .A(n954), .ZN(n1306) );
  AOI22_X1 U966 ( .A1(data_in[7]), .A2(n1650), .B1(n947), .B2(\mem[39][7] ), 
        .ZN(n954) );
  INV_X1 U967 ( .A(n1001), .ZN(n1265) );
  AOI22_X1 U968 ( .A1(data_in[0]), .A2(n1644), .B1(n1002), .B2(\mem[45][0] ), 
        .ZN(n1001) );
  INV_X1 U969 ( .A(n1003), .ZN(n1264) );
  AOI22_X1 U970 ( .A1(data_in[1]), .A2(n1644), .B1(n1002), .B2(\mem[45][1] ), 
        .ZN(n1003) );
  INV_X1 U971 ( .A(n1004), .ZN(n1263) );
  AOI22_X1 U972 ( .A1(data_in[2]), .A2(n1644), .B1(n1002), .B2(\mem[45][2] ), 
        .ZN(n1004) );
  INV_X1 U973 ( .A(n1005), .ZN(n1262) );
  AOI22_X1 U974 ( .A1(data_in[3]), .A2(n1644), .B1(n1002), .B2(\mem[45][3] ), 
        .ZN(n1005) );
  INV_X1 U975 ( .A(n1006), .ZN(n1261) );
  AOI22_X1 U976 ( .A1(data_in[4]), .A2(n1644), .B1(n1002), .B2(\mem[45][4] ), 
        .ZN(n1006) );
  INV_X1 U977 ( .A(n1007), .ZN(n1260) );
  AOI22_X1 U978 ( .A1(data_in[5]), .A2(n1644), .B1(n1002), .B2(\mem[45][5] ), 
        .ZN(n1007) );
  INV_X1 U979 ( .A(n1008), .ZN(n1259) );
  AOI22_X1 U980 ( .A1(data_in[6]), .A2(n1644), .B1(n1002), .B2(\mem[45][6] ), 
        .ZN(n1008) );
  INV_X1 U981 ( .A(n1009), .ZN(n1258) );
  AOI22_X1 U982 ( .A1(data_in[7]), .A2(n1644), .B1(n1002), .B2(\mem[45][7] ), 
        .ZN(n1009) );
  INV_X1 U983 ( .A(n1019), .ZN(n1249) );
  AOI22_X1 U984 ( .A1(data_in[0]), .A2(n1642), .B1(n1020), .B2(\mem[47][0] ), 
        .ZN(n1019) );
  INV_X1 U985 ( .A(n1021), .ZN(n1248) );
  AOI22_X1 U986 ( .A1(data_in[1]), .A2(n1642), .B1(n1020), .B2(\mem[47][1] ), 
        .ZN(n1021) );
  INV_X1 U987 ( .A(n1022), .ZN(n1247) );
  AOI22_X1 U988 ( .A1(data_in[2]), .A2(n1642), .B1(n1020), .B2(\mem[47][2] ), 
        .ZN(n1022) );
  INV_X1 U989 ( .A(n1023), .ZN(n1246) );
  AOI22_X1 U990 ( .A1(data_in[3]), .A2(n1642), .B1(n1020), .B2(\mem[47][3] ), 
        .ZN(n1023) );
  INV_X1 U991 ( .A(n1024), .ZN(n1245) );
  AOI22_X1 U992 ( .A1(data_in[4]), .A2(n1642), .B1(n1020), .B2(\mem[47][4] ), 
        .ZN(n1024) );
  INV_X1 U993 ( .A(n1025), .ZN(n1244) );
  AOI22_X1 U994 ( .A1(data_in[5]), .A2(n1642), .B1(n1020), .B2(\mem[47][5] ), 
        .ZN(n1025) );
  INV_X1 U995 ( .A(n1026), .ZN(n1243) );
  AOI22_X1 U996 ( .A1(data_in[6]), .A2(n1642), .B1(n1020), .B2(\mem[47][6] ), 
        .ZN(n1026) );
  INV_X1 U997 ( .A(n1027), .ZN(n1242) );
  AOI22_X1 U998 ( .A1(data_in[7]), .A2(n1642), .B1(n1020), .B2(\mem[47][7] ), 
        .ZN(n1027) );
  INV_X1 U999 ( .A(n1074), .ZN(n1201) );
  AOI22_X1 U1000 ( .A1(data_in[0]), .A2(n1636), .B1(n1075), .B2(\mem[53][0] ), 
        .ZN(n1074) );
  INV_X1 U1001 ( .A(n1076), .ZN(n1200) );
  AOI22_X1 U1002 ( .A1(data_in[1]), .A2(n1636), .B1(n1075), .B2(\mem[53][1] ), 
        .ZN(n1076) );
  INV_X1 U1003 ( .A(n1077), .ZN(n1199) );
  AOI22_X1 U1004 ( .A1(data_in[2]), .A2(n1636), .B1(n1075), .B2(\mem[53][2] ), 
        .ZN(n1077) );
  INV_X1 U1005 ( .A(n1078), .ZN(n1198) );
  AOI22_X1 U1006 ( .A1(data_in[3]), .A2(n1636), .B1(n1075), .B2(\mem[53][3] ), 
        .ZN(n1078) );
  INV_X1 U1007 ( .A(n1079), .ZN(n1197) );
  AOI22_X1 U1008 ( .A1(data_in[4]), .A2(n1636), .B1(n1075), .B2(\mem[53][4] ), 
        .ZN(n1079) );
  INV_X1 U1009 ( .A(n1080), .ZN(n1196) );
  AOI22_X1 U1010 ( .A1(data_in[5]), .A2(n1636), .B1(n1075), .B2(\mem[53][5] ), 
        .ZN(n1080) );
  INV_X1 U1011 ( .A(n1081), .ZN(n1195) );
  AOI22_X1 U1012 ( .A1(data_in[6]), .A2(n1636), .B1(n1075), .B2(\mem[53][6] ), 
        .ZN(n1081) );
  INV_X1 U1013 ( .A(n1082), .ZN(n1194) );
  AOI22_X1 U1014 ( .A1(data_in[7]), .A2(n1636), .B1(n1075), .B2(\mem[53][7] ), 
        .ZN(n1082) );
  INV_X1 U1015 ( .A(n1092), .ZN(n1185) );
  AOI22_X1 U1016 ( .A1(data_in[0]), .A2(n1634), .B1(n1093), .B2(\mem[55][0] ), 
        .ZN(n1092) );
  INV_X1 U1017 ( .A(n1094), .ZN(n1184) );
  AOI22_X1 U1018 ( .A1(data_in[1]), .A2(n1634), .B1(n1093), .B2(\mem[55][1] ), 
        .ZN(n1094) );
  INV_X1 U1019 ( .A(n1095), .ZN(n1183) );
  AOI22_X1 U1020 ( .A1(data_in[2]), .A2(n1634), .B1(n1093), .B2(\mem[55][2] ), 
        .ZN(n1095) );
  INV_X1 U1021 ( .A(n1096), .ZN(n1182) );
  AOI22_X1 U1022 ( .A1(data_in[3]), .A2(n1634), .B1(n1093), .B2(\mem[55][3] ), 
        .ZN(n1096) );
  INV_X1 U1023 ( .A(n1097), .ZN(n1181) );
  AOI22_X1 U1024 ( .A1(data_in[4]), .A2(n1634), .B1(n1093), .B2(\mem[55][4] ), 
        .ZN(n1097) );
  INV_X1 U1025 ( .A(n1098), .ZN(n1180) );
  AOI22_X1 U1026 ( .A1(data_in[5]), .A2(n1634), .B1(n1093), .B2(\mem[55][5] ), 
        .ZN(n1098) );
  INV_X1 U1027 ( .A(n1099), .ZN(n1179) );
  AOI22_X1 U1028 ( .A1(data_in[6]), .A2(n1634), .B1(n1093), .B2(\mem[55][6] ), 
        .ZN(n1099) );
  INV_X1 U1029 ( .A(n1100), .ZN(n1178) );
  AOI22_X1 U1030 ( .A1(data_in[7]), .A2(n1634), .B1(n1093), .B2(\mem[55][7] ), 
        .ZN(n1100) );
  INV_X1 U1031 ( .A(n1147), .ZN(n545) );
  AOI22_X1 U1032 ( .A1(data_in[0]), .A2(n1628), .B1(n1148), .B2(\mem[61][0] ), 
        .ZN(n1147) );
  INV_X1 U1033 ( .A(n1149), .ZN(n544) );
  AOI22_X1 U1034 ( .A1(data_in[1]), .A2(n1628), .B1(n1148), .B2(\mem[61][1] ), 
        .ZN(n1149) );
  INV_X1 U1035 ( .A(n1150), .ZN(n543) );
  AOI22_X1 U1036 ( .A1(data_in[2]), .A2(n1628), .B1(n1148), .B2(\mem[61][2] ), 
        .ZN(n1150) );
  INV_X1 U1037 ( .A(n1151), .ZN(n542) );
  AOI22_X1 U1038 ( .A1(data_in[3]), .A2(n1628), .B1(n1148), .B2(\mem[61][3] ), 
        .ZN(n1151) );
  INV_X1 U1039 ( .A(n1152), .ZN(n541) );
  AOI22_X1 U1040 ( .A1(data_in[4]), .A2(n1628), .B1(n1148), .B2(\mem[61][4] ), 
        .ZN(n1152) );
  INV_X1 U1041 ( .A(n1153), .ZN(n540) );
  AOI22_X1 U1042 ( .A1(data_in[5]), .A2(n1628), .B1(n1148), .B2(\mem[61][5] ), 
        .ZN(n1153) );
  INV_X1 U1043 ( .A(n1154), .ZN(n539) );
  AOI22_X1 U1044 ( .A1(data_in[6]), .A2(n1628), .B1(n1148), .B2(\mem[61][6] ), 
        .ZN(n1154) );
  INV_X1 U1045 ( .A(n1155), .ZN(n538) );
  AOI22_X1 U1046 ( .A1(data_in[7]), .A2(n1628), .B1(n1148), .B2(\mem[61][7] ), 
        .ZN(n1155) );
  INV_X1 U1047 ( .A(n1165), .ZN(n529) );
  AOI22_X1 U1048 ( .A1(data_in[0]), .A2(n1626), .B1(n1166), .B2(\mem[63][0] ), 
        .ZN(n1165) );
  INV_X1 U1049 ( .A(n1167), .ZN(n528) );
  AOI22_X1 U1050 ( .A1(data_in[1]), .A2(n1626), .B1(n1166), .B2(\mem[63][1] ), 
        .ZN(n1167) );
  INV_X1 U1051 ( .A(n1168), .ZN(n527) );
  AOI22_X1 U1052 ( .A1(data_in[2]), .A2(n1626), .B1(n1166), .B2(\mem[63][2] ), 
        .ZN(n1168) );
  INV_X1 U1053 ( .A(n1169), .ZN(n526) );
  AOI22_X1 U1054 ( .A1(data_in[3]), .A2(n1626), .B1(n1166), .B2(\mem[63][3] ), 
        .ZN(n1169) );
  INV_X1 U1055 ( .A(n1170), .ZN(n525) );
  AOI22_X1 U1056 ( .A1(data_in[4]), .A2(n1626), .B1(n1166), .B2(\mem[63][4] ), 
        .ZN(n1170) );
  INV_X1 U1057 ( .A(n1171), .ZN(n524) );
  AOI22_X1 U1058 ( .A1(data_in[5]), .A2(n1626), .B1(n1166), .B2(\mem[63][5] ), 
        .ZN(n1171) );
  INV_X1 U1059 ( .A(n1172), .ZN(n523) );
  AOI22_X1 U1060 ( .A1(data_in[6]), .A2(n1626), .B1(n1166), .B2(\mem[63][6] ), 
        .ZN(n1172) );
  INV_X1 U1061 ( .A(n1173), .ZN(n522) );
  AOI22_X1 U1062 ( .A1(data_in[7]), .A2(n1626), .B1(n1166), .B2(\mem[63][7] ), 
        .ZN(n1173) );
  INV_X1 U1063 ( .A(n582), .ZN(n1625) );
  AOI22_X1 U1064 ( .A1(n1689), .A2(data_in[0]), .B1(n583), .B2(\mem[0][0] ), 
        .ZN(n582) );
  INV_X1 U1065 ( .A(n584), .ZN(n1624) );
  AOI22_X1 U1066 ( .A1(n1689), .A2(data_in[1]), .B1(n583), .B2(\mem[0][1] ), 
        .ZN(n584) );
  INV_X1 U1067 ( .A(n585), .ZN(n1623) );
  AOI22_X1 U1068 ( .A1(n1689), .A2(data_in[2]), .B1(n583), .B2(\mem[0][2] ), 
        .ZN(n585) );
  INV_X1 U1069 ( .A(n586), .ZN(n1622) );
  AOI22_X1 U1070 ( .A1(n1689), .A2(data_in[3]), .B1(n583), .B2(\mem[0][3] ), 
        .ZN(n586) );
  INV_X1 U1071 ( .A(n587), .ZN(n1621) );
  AOI22_X1 U1072 ( .A1(n1689), .A2(data_in[4]), .B1(n583), .B2(\mem[0][4] ), 
        .ZN(n587) );
  INV_X1 U1073 ( .A(n588), .ZN(n1620) );
  AOI22_X1 U1074 ( .A1(n1689), .A2(data_in[5]), .B1(n583), .B2(\mem[0][5] ), 
        .ZN(n588) );
  INV_X1 U1075 ( .A(n589), .ZN(n1619) );
  AOI22_X1 U1076 ( .A1(n1689), .A2(data_in[6]), .B1(n583), .B2(\mem[0][6] ), 
        .ZN(n589) );
  INV_X1 U1077 ( .A(n590), .ZN(n1618) );
  AOI22_X1 U1078 ( .A1(n1689), .A2(data_in[7]), .B1(n583), .B2(\mem[0][7] ), 
        .ZN(n590) );
  INV_X1 U1079 ( .A(n593), .ZN(n1617) );
  AOI22_X1 U1080 ( .A1(data_in[0]), .A2(n1688), .B1(n594), .B2(\mem[1][0] ), 
        .ZN(n593) );
  INV_X1 U1081 ( .A(n595), .ZN(n1616) );
  AOI22_X1 U1082 ( .A1(data_in[1]), .A2(n1688), .B1(n594), .B2(\mem[1][1] ), 
        .ZN(n595) );
  INV_X1 U1083 ( .A(n596), .ZN(n1615) );
  AOI22_X1 U1084 ( .A1(data_in[2]), .A2(n1688), .B1(n594), .B2(\mem[1][2] ), 
        .ZN(n596) );
  INV_X1 U1085 ( .A(n597), .ZN(n1614) );
  AOI22_X1 U1086 ( .A1(data_in[3]), .A2(n1688), .B1(n594), .B2(\mem[1][3] ), 
        .ZN(n597) );
  INV_X1 U1087 ( .A(n598), .ZN(n1613) );
  AOI22_X1 U1088 ( .A1(data_in[4]), .A2(n1688), .B1(n594), .B2(\mem[1][4] ), 
        .ZN(n598) );
  INV_X1 U1089 ( .A(n599), .ZN(n1612) );
  AOI22_X1 U1090 ( .A1(data_in[5]), .A2(n1688), .B1(n594), .B2(\mem[1][5] ), 
        .ZN(n599) );
  INV_X1 U1091 ( .A(n600), .ZN(n1611) );
  AOI22_X1 U1092 ( .A1(data_in[6]), .A2(n1688), .B1(n594), .B2(\mem[1][6] ), 
        .ZN(n600) );
  INV_X1 U1093 ( .A(n601), .ZN(n1610) );
  AOI22_X1 U1094 ( .A1(data_in[7]), .A2(n1688), .B1(n594), .B2(\mem[1][7] ), 
        .ZN(n601) );
  INV_X1 U1095 ( .A(n603), .ZN(n1609) );
  AOI22_X1 U1096 ( .A1(data_in[0]), .A2(n1687), .B1(n604), .B2(\mem[2][0] ), 
        .ZN(n603) );
  INV_X1 U1097 ( .A(n605), .ZN(n1608) );
  AOI22_X1 U1098 ( .A1(data_in[1]), .A2(n1687), .B1(n604), .B2(\mem[2][1] ), 
        .ZN(n605) );
  INV_X1 U1099 ( .A(n606), .ZN(n1607) );
  AOI22_X1 U1100 ( .A1(data_in[2]), .A2(n1687), .B1(n604), .B2(\mem[2][2] ), 
        .ZN(n606) );
  INV_X1 U1101 ( .A(n607), .ZN(n1606) );
  AOI22_X1 U1102 ( .A1(data_in[3]), .A2(n1687), .B1(n604), .B2(\mem[2][3] ), 
        .ZN(n607) );
  INV_X1 U1103 ( .A(n608), .ZN(n1605) );
  AOI22_X1 U1104 ( .A1(data_in[4]), .A2(n1687), .B1(n604), .B2(\mem[2][4] ), 
        .ZN(n608) );
  INV_X1 U1105 ( .A(n609), .ZN(n1604) );
  AOI22_X1 U1106 ( .A1(data_in[5]), .A2(n1687), .B1(n604), .B2(\mem[2][5] ), 
        .ZN(n609) );
  INV_X1 U1107 ( .A(n610), .ZN(n1603) );
  AOI22_X1 U1108 ( .A1(data_in[6]), .A2(n1687), .B1(n604), .B2(\mem[2][6] ), 
        .ZN(n610) );
  INV_X1 U1109 ( .A(n611), .ZN(n1602) );
  AOI22_X1 U1110 ( .A1(data_in[7]), .A2(n1687), .B1(n604), .B2(\mem[2][7] ), 
        .ZN(n611) );
  INV_X1 U1111 ( .A(n613), .ZN(n1601) );
  AOI22_X1 U1112 ( .A1(data_in[0]), .A2(n1686), .B1(n614), .B2(\mem[3][0] ), 
        .ZN(n613) );
  INV_X1 U1113 ( .A(n615), .ZN(n1600) );
  AOI22_X1 U1114 ( .A1(data_in[1]), .A2(n1686), .B1(n614), .B2(\mem[3][1] ), 
        .ZN(n615) );
  INV_X1 U1115 ( .A(n616), .ZN(n1599) );
  AOI22_X1 U1116 ( .A1(data_in[2]), .A2(n1686), .B1(n614), .B2(\mem[3][2] ), 
        .ZN(n616) );
  INV_X1 U1117 ( .A(n617), .ZN(n1598) );
  AOI22_X1 U1118 ( .A1(data_in[3]), .A2(n1686), .B1(n614), .B2(\mem[3][3] ), 
        .ZN(n617) );
  INV_X1 U1119 ( .A(n618), .ZN(n1597) );
  AOI22_X1 U1120 ( .A1(data_in[4]), .A2(n1686), .B1(n614), .B2(\mem[3][4] ), 
        .ZN(n618) );
  INV_X1 U1121 ( .A(n619), .ZN(n1596) );
  AOI22_X1 U1122 ( .A1(data_in[5]), .A2(n1686), .B1(n614), .B2(\mem[3][5] ), 
        .ZN(n619) );
  INV_X1 U1123 ( .A(n620), .ZN(n1595) );
  AOI22_X1 U1124 ( .A1(data_in[6]), .A2(n1686), .B1(n614), .B2(\mem[3][6] ), 
        .ZN(n620) );
  INV_X1 U1125 ( .A(n621), .ZN(n1594) );
  AOI22_X1 U1126 ( .A1(data_in[7]), .A2(n1686), .B1(n614), .B2(\mem[3][7] ), 
        .ZN(n621) );
  INV_X1 U1127 ( .A(n623), .ZN(n1593) );
  AOI22_X1 U1128 ( .A1(data_in[0]), .A2(n1685), .B1(n624), .B2(\mem[4][0] ), 
        .ZN(n623) );
  INV_X1 U1129 ( .A(n625), .ZN(n1592) );
  AOI22_X1 U1130 ( .A1(data_in[1]), .A2(n1685), .B1(n624), .B2(\mem[4][1] ), 
        .ZN(n625) );
  INV_X1 U1131 ( .A(n626), .ZN(n1591) );
  AOI22_X1 U1132 ( .A1(data_in[2]), .A2(n1685), .B1(n624), .B2(\mem[4][2] ), 
        .ZN(n626) );
  INV_X1 U1133 ( .A(n627), .ZN(n1590) );
  AOI22_X1 U1134 ( .A1(data_in[3]), .A2(n1685), .B1(n624), .B2(\mem[4][3] ), 
        .ZN(n627) );
  INV_X1 U1135 ( .A(n628), .ZN(n1589) );
  AOI22_X1 U1136 ( .A1(data_in[4]), .A2(n1685), .B1(n624), .B2(\mem[4][4] ), 
        .ZN(n628) );
  INV_X1 U1137 ( .A(n629), .ZN(n1588) );
  AOI22_X1 U1138 ( .A1(data_in[5]), .A2(n1685), .B1(n624), .B2(\mem[4][5] ), 
        .ZN(n629) );
  INV_X1 U1139 ( .A(n630), .ZN(n1587) );
  AOI22_X1 U1140 ( .A1(data_in[6]), .A2(n1685), .B1(n624), .B2(\mem[4][6] ), 
        .ZN(n630) );
  INV_X1 U1141 ( .A(n631), .ZN(n1586) );
  AOI22_X1 U1142 ( .A1(data_in[7]), .A2(n1685), .B1(n624), .B2(\mem[4][7] ), 
        .ZN(n631) );
  INV_X1 U1143 ( .A(n633), .ZN(n1585) );
  AOI22_X1 U1144 ( .A1(data_in[0]), .A2(n1684), .B1(n634), .B2(\mem[5][0] ), 
        .ZN(n633) );
  INV_X1 U1145 ( .A(n635), .ZN(n1584) );
  AOI22_X1 U1146 ( .A1(data_in[1]), .A2(n1684), .B1(n634), .B2(\mem[5][1] ), 
        .ZN(n635) );
  INV_X1 U1147 ( .A(n636), .ZN(n1583) );
  AOI22_X1 U1148 ( .A1(data_in[2]), .A2(n1684), .B1(n634), .B2(\mem[5][2] ), 
        .ZN(n636) );
  INV_X1 U1149 ( .A(n637), .ZN(n1582) );
  AOI22_X1 U1150 ( .A1(data_in[3]), .A2(n1684), .B1(n634), .B2(\mem[5][3] ), 
        .ZN(n637) );
  INV_X1 U1151 ( .A(n638), .ZN(n1581) );
  AOI22_X1 U1152 ( .A1(data_in[4]), .A2(n1684), .B1(n634), .B2(\mem[5][4] ), 
        .ZN(n638) );
  INV_X1 U1153 ( .A(n639), .ZN(n1580) );
  AOI22_X1 U1154 ( .A1(data_in[5]), .A2(n1684), .B1(n634), .B2(\mem[5][5] ), 
        .ZN(n639) );
  INV_X1 U1155 ( .A(n640), .ZN(n1579) );
  AOI22_X1 U1156 ( .A1(data_in[6]), .A2(n1684), .B1(n634), .B2(\mem[5][6] ), 
        .ZN(n640) );
  INV_X1 U1157 ( .A(n641), .ZN(n1578) );
  AOI22_X1 U1158 ( .A1(data_in[7]), .A2(n1684), .B1(n634), .B2(\mem[5][7] ), 
        .ZN(n641) );
  INV_X1 U1159 ( .A(n643), .ZN(n1577) );
  AOI22_X1 U1160 ( .A1(data_in[0]), .A2(n1683), .B1(n644), .B2(\mem[6][0] ), 
        .ZN(n643) );
  INV_X1 U1161 ( .A(n645), .ZN(n1576) );
  AOI22_X1 U1162 ( .A1(data_in[1]), .A2(n1683), .B1(n644), .B2(\mem[6][1] ), 
        .ZN(n645) );
  INV_X1 U1163 ( .A(n646), .ZN(n1575) );
  AOI22_X1 U1164 ( .A1(data_in[2]), .A2(n1683), .B1(n644), .B2(\mem[6][2] ), 
        .ZN(n646) );
  INV_X1 U1165 ( .A(n647), .ZN(n1574) );
  AOI22_X1 U1166 ( .A1(data_in[3]), .A2(n1683), .B1(n644), .B2(\mem[6][3] ), 
        .ZN(n647) );
  INV_X1 U1167 ( .A(n648), .ZN(n1573) );
  AOI22_X1 U1168 ( .A1(data_in[4]), .A2(n1683), .B1(n644), .B2(\mem[6][4] ), 
        .ZN(n648) );
  INV_X1 U1169 ( .A(n649), .ZN(n1572) );
  AOI22_X1 U1170 ( .A1(data_in[5]), .A2(n1683), .B1(n644), .B2(\mem[6][5] ), 
        .ZN(n649) );
  INV_X1 U1171 ( .A(n650), .ZN(n1571) );
  AOI22_X1 U1172 ( .A1(data_in[6]), .A2(n1683), .B1(n644), .B2(\mem[6][6] ), 
        .ZN(n650) );
  INV_X1 U1173 ( .A(n651), .ZN(n1570) );
  AOI22_X1 U1174 ( .A1(data_in[7]), .A2(n1683), .B1(n644), .B2(\mem[6][7] ), 
        .ZN(n651) );
  INV_X1 U1175 ( .A(n653), .ZN(n1569) );
  AOI22_X1 U1176 ( .A1(data_in[0]), .A2(n1682), .B1(n654), .B2(\mem[7][0] ), 
        .ZN(n653) );
  INV_X1 U1177 ( .A(n655), .ZN(n1568) );
  AOI22_X1 U1178 ( .A1(data_in[1]), .A2(n1682), .B1(n654), .B2(\mem[7][1] ), 
        .ZN(n655) );
  INV_X1 U1179 ( .A(n656), .ZN(n1567) );
  AOI22_X1 U1180 ( .A1(data_in[2]), .A2(n1682), .B1(n654), .B2(\mem[7][2] ), 
        .ZN(n656) );
  INV_X1 U1181 ( .A(n657), .ZN(n1566) );
  AOI22_X1 U1182 ( .A1(data_in[3]), .A2(n1682), .B1(n654), .B2(\mem[7][3] ), 
        .ZN(n657) );
  INV_X1 U1183 ( .A(n658), .ZN(n1565) );
  AOI22_X1 U1184 ( .A1(data_in[4]), .A2(n1682), .B1(n654), .B2(\mem[7][4] ), 
        .ZN(n658) );
  INV_X1 U1185 ( .A(n659), .ZN(n1564) );
  AOI22_X1 U1186 ( .A1(data_in[5]), .A2(n1682), .B1(n654), .B2(\mem[7][5] ), 
        .ZN(n659) );
  INV_X1 U1187 ( .A(n660), .ZN(n1563) );
  AOI22_X1 U1188 ( .A1(data_in[6]), .A2(n1682), .B1(n654), .B2(\mem[7][6] ), 
        .ZN(n660) );
  INV_X1 U1189 ( .A(n661), .ZN(n1562) );
  AOI22_X1 U1190 ( .A1(data_in[7]), .A2(n1682), .B1(n654), .B2(\mem[7][7] ), 
        .ZN(n661) );
  MUX2_X1 U1191 ( .A(\mem[62][0] ), .B(\mem[63][0] ), .S(n511), .Z(n3) );
  MUX2_X1 U1192 ( .A(\mem[60][0] ), .B(\mem[61][0] ), .S(n511), .Z(n4) );
  MUX2_X1 U1193 ( .A(n4), .B(n3), .S(n503), .Z(n5) );
  MUX2_X1 U1194 ( .A(\mem[58][0] ), .B(\mem[59][0] ), .S(n511), .Z(n6) );
  MUX2_X1 U1195 ( .A(\mem[56][0] ), .B(\mem[57][0] ), .S(n513), .Z(n7) );
  MUX2_X1 U1196 ( .A(n7), .B(n6), .S(n503), .Z(n8) );
  MUX2_X1 U1197 ( .A(n8), .B(n5), .S(n502), .Z(n9) );
  MUX2_X1 U1198 ( .A(\mem[54][0] ), .B(\mem[55][0] ), .S(n511), .Z(n10) );
  MUX2_X1 U1199 ( .A(\mem[52][0] ), .B(\mem[53][0] ), .S(n511), .Z(n11) );
  MUX2_X1 U1200 ( .A(n11), .B(n10), .S(n503), .Z(n12) );
  MUX2_X1 U1201 ( .A(\mem[50][0] ), .B(\mem[51][0] ), .S(n510), .Z(n13) );
  MUX2_X1 U1202 ( .A(\mem[48][0] ), .B(\mem[49][0] ), .S(n510), .Z(n14) );
  MUX2_X1 U1203 ( .A(n14), .B(n13), .S(n503), .Z(n15) );
  MUX2_X1 U1204 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U1205 ( .A(n16), .B(n9), .S(n499), .Z(n17) );
  MUX2_X1 U1206 ( .A(\mem[46][0] ), .B(\mem[47][0] ), .S(n511), .Z(n18) );
  MUX2_X1 U1207 ( .A(\mem[44][0] ), .B(\mem[45][0] ), .S(n511), .Z(n19) );
  MUX2_X1 U1208 ( .A(n19), .B(n18), .S(n503), .Z(n20) );
  MUX2_X1 U1209 ( .A(\mem[42][0] ), .B(\mem[43][0] ), .S(n510), .Z(n21) );
  MUX2_X1 U1210 ( .A(\mem[40][0] ), .B(\mem[41][0] ), .S(n513), .Z(n22) );
  MUX2_X1 U1211 ( .A(n22), .B(n21), .S(n503), .Z(n23) );
  MUX2_X1 U1212 ( .A(n23), .B(n20), .S(n501), .Z(n24) );
  MUX2_X1 U1213 ( .A(\mem[38][0] ), .B(\mem[39][0] ), .S(n510), .Z(n25) );
  MUX2_X1 U1214 ( .A(\mem[36][0] ), .B(\mem[37][0] ), .S(n510), .Z(n26) );
  MUX2_X1 U1215 ( .A(n26), .B(n25), .S(n503), .Z(n27) );
  MUX2_X1 U1216 ( .A(\mem[34][0] ), .B(\mem[35][0] ), .S(n510), .Z(n28) );
  MUX2_X1 U1217 ( .A(\mem[32][0] ), .B(\mem[33][0] ), .S(n510), .Z(n29) );
  MUX2_X1 U1218 ( .A(n29), .B(n28), .S(n503), .Z(n30) );
  MUX2_X1 U1219 ( .A(n30), .B(n27), .S(N12), .Z(n31) );
  MUX2_X1 U1220 ( .A(n31), .B(n24), .S(n499), .Z(n32) );
  MUX2_X1 U1221 ( .A(n32), .B(n17), .S(N14), .Z(n33) );
  MUX2_X1 U1222 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n510), .Z(n34) );
  MUX2_X1 U1223 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n510), .Z(n35) );
  MUX2_X1 U1224 ( .A(n35), .B(n34), .S(n504), .Z(n36) );
  MUX2_X1 U1225 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n510), .Z(n37) );
  MUX2_X1 U1226 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n510), .Z(n38) );
  MUX2_X1 U1227 ( .A(n38), .B(n37), .S(n504), .Z(n39) );
  MUX2_X1 U1228 ( .A(n39), .B(n36), .S(n500), .Z(n40) );
  MUX2_X1 U1229 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n510), .Z(n41) );
  MUX2_X1 U1230 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n510), .Z(n42) );
  MUX2_X1 U1231 ( .A(n42), .B(n41), .S(n504), .Z(n43) );
  MUX2_X1 U1232 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n510), .Z(n44) );
  MUX2_X1 U1233 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n510), .Z(n45) );
  MUX2_X1 U1234 ( .A(n45), .B(n44), .S(n504), .Z(n46) );
  MUX2_X1 U1235 ( .A(n46), .B(n43), .S(N12), .Z(n47) );
  MUX2_X1 U1236 ( .A(n47), .B(n40), .S(n499), .Z(n48) );
  MUX2_X1 U1237 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n510), .Z(n49) );
  MUX2_X1 U1238 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n510), .Z(n50) );
  MUX2_X1 U1239 ( .A(n50), .B(n49), .S(n504), .Z(n51) );
  MUX2_X1 U1240 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n510), .Z(n52) );
  MUX2_X1 U1241 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n510), .Z(n53) );
  MUX2_X1 U1242 ( .A(n53), .B(n52), .S(n504), .Z(n54) );
  MUX2_X1 U1243 ( .A(n54), .B(n51), .S(n500), .Z(n55) );
  MUX2_X1 U1244 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n513), .Z(n56) );
  MUX2_X1 U1245 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n511), .Z(n57) );
  MUX2_X1 U1246 ( .A(n57), .B(n56), .S(n504), .Z(n58) );
  MUX2_X1 U1247 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n512), .Z(n59) );
  MUX2_X1 U1248 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n513), .Z(n60) );
  MUX2_X1 U1249 ( .A(n60), .B(n59), .S(n504), .Z(n61) );
  MUX2_X1 U1250 ( .A(n61), .B(n58), .S(N12), .Z(n62) );
  MUX2_X1 U1251 ( .A(n62), .B(n55), .S(n499), .Z(n63) );
  MUX2_X1 U1252 ( .A(n63), .B(n48), .S(N14), .Z(n64) );
  MUX2_X1 U1253 ( .A(n64), .B(n33), .S(N15), .Z(N23) );
  MUX2_X1 U1254 ( .A(\mem[62][1] ), .B(\mem[63][1] ), .S(n513), .Z(n65) );
  MUX2_X1 U1255 ( .A(\mem[60][1] ), .B(\mem[61][1] ), .S(n512), .Z(n66) );
  MUX2_X1 U1256 ( .A(n66), .B(n65), .S(n504), .Z(n67) );
  MUX2_X1 U1257 ( .A(\mem[58][1] ), .B(\mem[59][1] ), .S(n511), .Z(n68) );
  MUX2_X1 U1258 ( .A(\mem[56][1] ), .B(\mem[57][1] ), .S(n511), .Z(n69) );
  MUX2_X1 U1259 ( .A(n69), .B(n68), .S(n504), .Z(n70) );
  MUX2_X1 U1260 ( .A(n70), .B(n67), .S(N12), .Z(n71) );
  MUX2_X1 U1261 ( .A(\mem[54][1] ), .B(\mem[55][1] ), .S(n516), .Z(n72) );
  MUX2_X1 U1262 ( .A(\mem[52][1] ), .B(\mem[53][1] ), .S(n513), .Z(n73) );
  MUX2_X1 U1263 ( .A(n73), .B(n72), .S(n504), .Z(n74) );
  MUX2_X1 U1264 ( .A(\mem[50][1] ), .B(\mem[51][1] ), .S(n511), .Z(n75) );
  MUX2_X1 U1265 ( .A(\mem[48][1] ), .B(\mem[49][1] ), .S(n512), .Z(n76) );
  MUX2_X1 U1266 ( .A(n76), .B(n75), .S(n504), .Z(n77) );
  MUX2_X1 U1267 ( .A(n77), .B(n74), .S(n502), .Z(n78) );
  MUX2_X1 U1268 ( .A(n78), .B(n71), .S(n499), .Z(n79) );
  MUX2_X1 U1269 ( .A(\mem[46][1] ), .B(\mem[47][1] ), .S(n510), .Z(n80) );
  MUX2_X1 U1270 ( .A(\mem[44][1] ), .B(\mem[45][1] ), .S(n513), .Z(n81) );
  MUX2_X1 U1271 ( .A(n81), .B(n80), .S(n508), .Z(n82) );
  MUX2_X1 U1272 ( .A(\mem[42][1] ), .B(\mem[43][1] ), .S(n514), .Z(n83) );
  MUX2_X1 U1273 ( .A(\mem[40][1] ), .B(\mem[41][1] ), .S(n512), .Z(n84) );
  MUX2_X1 U1274 ( .A(n84), .B(n83), .S(N11), .Z(n85) );
  MUX2_X1 U1275 ( .A(n85), .B(n82), .S(n501), .Z(n86) );
  MUX2_X1 U1276 ( .A(\mem[38][1] ), .B(\mem[39][1] ), .S(n510), .Z(n87) );
  MUX2_X1 U1277 ( .A(\mem[36][1] ), .B(\mem[37][1] ), .S(n511), .Z(n88) );
  MUX2_X1 U1278 ( .A(n88), .B(n87), .S(n509), .Z(n89) );
  MUX2_X1 U1279 ( .A(\mem[34][1] ), .B(\mem[35][1] ), .S(n510), .Z(n90) );
  MUX2_X1 U1280 ( .A(\mem[32][1] ), .B(\mem[33][1] ), .S(n510), .Z(n91) );
  MUX2_X1 U1281 ( .A(n91), .B(n90), .S(N11), .Z(n92) );
  MUX2_X1 U1282 ( .A(n92), .B(n89), .S(n500), .Z(n93) );
  MUX2_X1 U1283 ( .A(n93), .B(n86), .S(n499), .Z(n94) );
  MUX2_X1 U1284 ( .A(n94), .B(n79), .S(N14), .Z(n95) );
  MUX2_X1 U1285 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n513), .Z(n96) );
  MUX2_X1 U1286 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n513), .Z(n97) );
  MUX2_X1 U1287 ( .A(n97), .B(n96), .S(n508), .Z(n98) );
  MUX2_X1 U1288 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n512), .Z(n99) );
  MUX2_X1 U1289 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n511), .Z(n100) );
  MUX2_X1 U1290 ( .A(n100), .B(n99), .S(N11), .Z(n101) );
  MUX2_X1 U1291 ( .A(n101), .B(n98), .S(N12), .Z(n102) );
  MUX2_X1 U1292 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n511), .Z(n103) );
  MUX2_X1 U1293 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n512), .Z(n104) );
  MUX2_X1 U1294 ( .A(n104), .B(n103), .S(n508), .Z(n105) );
  MUX2_X1 U1295 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n510), .Z(n106) );
  MUX2_X1 U1296 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n513), .Z(n107) );
  MUX2_X1 U1297 ( .A(n107), .B(n106), .S(N11), .Z(n108) );
  MUX2_X1 U1298 ( .A(n108), .B(n105), .S(N12), .Z(n109) );
  MUX2_X1 U1299 ( .A(n109), .B(n102), .S(n499), .Z(n110) );
  MUX2_X1 U1300 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n513), .Z(n111) );
  MUX2_X1 U1301 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n513), .Z(n112) );
  MUX2_X1 U1302 ( .A(n112), .B(n111), .S(n503), .Z(n113) );
  MUX2_X1 U1303 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n513), .Z(n114) );
  MUX2_X1 U1304 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n512), .Z(n115) );
  MUX2_X1 U1305 ( .A(n115), .B(n114), .S(n506), .Z(n116) );
  MUX2_X1 U1306 ( .A(n116), .B(n113), .S(N12), .Z(n117) );
  MUX2_X1 U1307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n510), .Z(n118) );
  MUX2_X1 U1308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n516), .Z(n119) );
  MUX2_X1 U1309 ( .A(n119), .B(n118), .S(N11), .Z(n120) );
  MUX2_X1 U1310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n121) );
  MUX2_X1 U1311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n512), .Z(n122) );
  MUX2_X1 U1312 ( .A(n122), .B(n121), .S(N11), .Z(n123) );
  MUX2_X1 U1313 ( .A(n123), .B(n120), .S(N12), .Z(n124) );
  MUX2_X1 U1314 ( .A(n124), .B(n117), .S(n499), .Z(n125) );
  MUX2_X1 U1315 ( .A(n125), .B(n110), .S(N14), .Z(n126) );
  MUX2_X1 U1316 ( .A(\mem[62][2] ), .B(\mem[63][2] ), .S(n510), .Z(n127) );
  MUX2_X1 U1317 ( .A(\mem[60][2] ), .B(\mem[61][2] ), .S(n512), .Z(n128) );
  MUX2_X1 U1318 ( .A(n128), .B(n127), .S(n505), .Z(n129) );
  MUX2_X1 U1319 ( .A(\mem[58][2] ), .B(\mem[59][2] ), .S(n511), .Z(n130) );
  MUX2_X1 U1320 ( .A(\mem[56][2] ), .B(\mem[57][2] ), .S(n510), .Z(n131) );
  MUX2_X1 U1321 ( .A(n131), .B(n130), .S(n505), .Z(n132) );
  MUX2_X1 U1322 ( .A(n132), .B(n129), .S(n502), .Z(n133) );
  MUX2_X1 U1323 ( .A(\mem[54][2] ), .B(\mem[55][2] ), .S(n516), .Z(n134) );
  MUX2_X1 U1324 ( .A(\mem[52][2] ), .B(\mem[53][2] ), .S(n511), .Z(n135) );
  MUX2_X1 U1325 ( .A(n135), .B(n134), .S(n505), .Z(n136) );
  MUX2_X1 U1326 ( .A(\mem[50][2] ), .B(\mem[51][2] ), .S(n512), .Z(n137) );
  MUX2_X1 U1327 ( .A(\mem[48][2] ), .B(\mem[49][2] ), .S(N10), .Z(n138) );
  MUX2_X1 U1328 ( .A(n138), .B(n137), .S(n505), .Z(n139) );
  MUX2_X1 U1329 ( .A(n139), .B(n136), .S(n501), .Z(n140) );
  MUX2_X1 U1330 ( .A(n140), .B(n133), .S(n499), .Z(n141) );
  MUX2_X1 U1331 ( .A(\mem[46][2] ), .B(\mem[47][2] ), .S(n510), .Z(n142) );
  MUX2_X1 U1332 ( .A(\mem[44][2] ), .B(\mem[45][2] ), .S(n511), .Z(n143) );
  MUX2_X1 U1333 ( .A(n143), .B(n142), .S(n505), .Z(n144) );
  MUX2_X1 U1334 ( .A(\mem[42][2] ), .B(\mem[43][2] ), .S(n510), .Z(n145) );
  MUX2_X1 U1335 ( .A(\mem[40][2] ), .B(\mem[41][2] ), .S(n511), .Z(n146) );
  MUX2_X1 U1336 ( .A(n146), .B(n145), .S(n505), .Z(n147) );
  MUX2_X1 U1337 ( .A(n147), .B(n144), .S(n500), .Z(n148) );
  MUX2_X1 U1338 ( .A(\mem[38][2] ), .B(\mem[39][2] ), .S(n510), .Z(n149) );
  MUX2_X1 U1339 ( .A(\mem[36][2] ), .B(\mem[37][2] ), .S(n511), .Z(n150) );
  MUX2_X1 U1340 ( .A(n150), .B(n149), .S(n505), .Z(n151) );
  MUX2_X1 U1341 ( .A(\mem[34][2] ), .B(\mem[35][2] ), .S(n512), .Z(n152) );
  MUX2_X1 U1342 ( .A(\mem[32][2] ), .B(\mem[33][2] ), .S(n513), .Z(n153) );
  MUX2_X1 U1343 ( .A(n153), .B(n152), .S(n505), .Z(n154) );
  MUX2_X1 U1344 ( .A(n154), .B(n151), .S(n502), .Z(n155) );
  MUX2_X1 U1345 ( .A(n155), .B(n148), .S(N13), .Z(n156) );
  MUX2_X1 U1346 ( .A(n156), .B(n141), .S(N14), .Z(n157) );
  MUX2_X1 U1347 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n510), .Z(n158) );
  MUX2_X1 U1348 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(N10), .Z(n159) );
  MUX2_X1 U1349 ( .A(n159), .B(n158), .S(n505), .Z(n160) );
  MUX2_X1 U1350 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n511), .Z(n161) );
  MUX2_X1 U1351 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n511), .Z(n162) );
  MUX2_X1 U1352 ( .A(n162), .B(n161), .S(n505), .Z(n163) );
  MUX2_X1 U1353 ( .A(n163), .B(n160), .S(n501), .Z(n164) );
  MUX2_X1 U1354 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n510), .Z(n165) );
  MUX2_X1 U1355 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n511), .Z(n166) );
  MUX2_X1 U1356 ( .A(n166), .B(n165), .S(n505), .Z(n167) );
  MUX2_X1 U1357 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n516), .Z(n168) );
  MUX2_X1 U1358 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n513), .Z(n169) );
  MUX2_X1 U1359 ( .A(n169), .B(n168), .S(n505), .Z(n170) );
  MUX2_X1 U1360 ( .A(n170), .B(n167), .S(n501), .Z(n171) );
  MUX2_X1 U1361 ( .A(n171), .B(n164), .S(N13), .Z(n172) );
  MUX2_X1 U1362 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n511), .Z(n173) );
  MUX2_X1 U1363 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n511), .Z(n174) );
  MUX2_X1 U1364 ( .A(n174), .B(n173), .S(n503), .Z(n175) );
  MUX2_X1 U1365 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n512), .Z(n176) );
  MUX2_X1 U1366 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n177) );
  MUX2_X1 U1367 ( .A(n177), .B(n176), .S(n503), .Z(n178) );
  MUX2_X1 U1368 ( .A(n178), .B(n175), .S(n502), .Z(n179) );
  MUX2_X1 U1369 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n512), .Z(n180) );
  MUX2_X1 U1370 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n510), .Z(n181) );
  MUX2_X1 U1371 ( .A(n181), .B(n180), .S(n503), .Z(n182) );
  MUX2_X1 U1372 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n513), .Z(n183) );
  MUX2_X1 U1373 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n511), .Z(n184) );
  MUX2_X1 U1374 ( .A(n184), .B(n183), .S(N11), .Z(n185) );
  MUX2_X1 U1375 ( .A(n185), .B(n182), .S(n500), .Z(n186) );
  MUX2_X1 U1376 ( .A(n186), .B(n179), .S(N13), .Z(n187) );
  MUX2_X1 U1377 ( .A(n187), .B(n172), .S(N14), .Z(n188) );
  MUX2_X1 U1378 ( .A(n188), .B(n157), .S(N15), .Z(N21) );
  MUX2_X1 U1379 ( .A(\mem[62][3] ), .B(\mem[63][3] ), .S(N10), .Z(n189) );
  MUX2_X1 U1380 ( .A(\mem[60][3] ), .B(\mem[61][3] ), .S(n513), .Z(n190) );
  MUX2_X1 U1381 ( .A(n190), .B(n189), .S(n507), .Z(n191) );
  MUX2_X1 U1382 ( .A(\mem[58][3] ), .B(\mem[59][3] ), .S(n510), .Z(n192) );
  MUX2_X1 U1383 ( .A(\mem[56][3] ), .B(\mem[57][3] ), .S(n513), .Z(n193) );
  MUX2_X1 U1384 ( .A(n193), .B(n192), .S(n508), .Z(n194) );
  MUX2_X1 U1385 ( .A(n194), .B(n191), .S(n501), .Z(n195) );
  MUX2_X1 U1386 ( .A(\mem[54][3] ), .B(\mem[55][3] ), .S(n513), .Z(n196) );
  MUX2_X1 U1387 ( .A(\mem[52][3] ), .B(\mem[53][3] ), .S(n511), .Z(n197) );
  MUX2_X1 U1388 ( .A(n197), .B(n196), .S(n506), .Z(n198) );
  MUX2_X1 U1389 ( .A(\mem[50][3] ), .B(\mem[51][3] ), .S(N10), .Z(n199) );
  MUX2_X1 U1390 ( .A(\mem[48][3] ), .B(\mem[49][3] ), .S(n510), .Z(n200) );
  MUX2_X1 U1391 ( .A(n200), .B(n199), .S(N11), .Z(n201) );
  MUX2_X1 U1392 ( .A(n201), .B(n198), .S(n500), .Z(n202) );
  MUX2_X1 U1393 ( .A(n202), .B(n195), .S(N13), .Z(n203) );
  MUX2_X1 U1394 ( .A(\mem[46][3] ), .B(\mem[47][3] ), .S(n511), .Z(n204) );
  MUX2_X1 U1395 ( .A(\mem[44][3] ), .B(\mem[45][3] ), .S(n513), .Z(n205) );
  MUX2_X1 U1396 ( .A(n205), .B(n204), .S(n507), .Z(n206) );
  MUX2_X1 U1397 ( .A(\mem[42][3] ), .B(\mem[43][3] ), .S(n511), .Z(n207) );
  MUX2_X1 U1398 ( .A(\mem[40][3] ), .B(\mem[41][3] ), .S(n511), .Z(n208) );
  MUX2_X1 U1399 ( .A(n208), .B(n207), .S(n506), .Z(n209) );
  MUX2_X1 U1400 ( .A(n209), .B(n206), .S(n502), .Z(n210) );
  MUX2_X1 U1401 ( .A(\mem[38][3] ), .B(\mem[39][3] ), .S(n511), .Z(n211) );
  MUX2_X1 U1402 ( .A(\mem[36][3] ), .B(\mem[37][3] ), .S(n516), .Z(n212) );
  MUX2_X1 U1403 ( .A(n212), .B(n211), .S(n509), .Z(n213) );
  MUX2_X1 U1404 ( .A(\mem[34][3] ), .B(\mem[35][3] ), .S(n513), .Z(n214) );
  MUX2_X1 U1405 ( .A(\mem[32][3] ), .B(\mem[33][3] ), .S(N10), .Z(n215) );
  MUX2_X1 U1406 ( .A(n215), .B(n214), .S(n507), .Z(n216) );
  MUX2_X1 U1407 ( .A(n216), .B(n213), .S(n501), .Z(n217) );
  MUX2_X1 U1408 ( .A(n217), .B(n210), .S(N13), .Z(n218) );
  MUX2_X1 U1409 ( .A(n218), .B(n203), .S(N14), .Z(n219) );
  MUX2_X1 U1410 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n513), .Z(n220) );
  MUX2_X1 U1411 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n512), .Z(n221) );
  MUX2_X1 U1412 ( .A(n221), .B(n220), .S(n503), .Z(n222) );
  MUX2_X1 U1413 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n512), .Z(n223) );
  MUX2_X1 U1414 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n511), .Z(n224) );
  MUX2_X1 U1415 ( .A(n224), .B(n223), .S(n504), .Z(n225) );
  MUX2_X1 U1416 ( .A(n225), .B(n222), .S(n500), .Z(n226) );
  MUX2_X1 U1417 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n510), .Z(n227) );
  MUX2_X1 U1418 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n510), .Z(n228) );
  MUX2_X1 U1419 ( .A(n228), .B(n227), .S(n504), .Z(n229) );
  MUX2_X1 U1420 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n511), .Z(n230) );
  MUX2_X1 U1421 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n511), .Z(n231) );
  MUX2_X1 U1422 ( .A(n231), .B(n230), .S(n503), .Z(n232) );
  MUX2_X1 U1423 ( .A(n232), .B(n229), .S(n500), .Z(n233) );
  MUX2_X1 U1424 ( .A(n233), .B(n226), .S(N13), .Z(n234) );
  MUX2_X1 U1425 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n512), .Z(n235) );
  MUX2_X1 U1426 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n516), .Z(n236) );
  MUX2_X1 U1427 ( .A(n236), .B(n235), .S(n503), .Z(n237) );
  MUX2_X1 U1428 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n512), .Z(n238) );
  MUX2_X1 U1429 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n511), .Z(n239) );
  MUX2_X1 U1430 ( .A(n239), .B(n238), .S(n504), .Z(n240) );
  MUX2_X1 U1431 ( .A(n240), .B(n237), .S(n500), .Z(n241) );
  MUX2_X1 U1432 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n513), .Z(n242) );
  MUX2_X1 U1433 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n512), .Z(n243) );
  MUX2_X1 U1434 ( .A(n243), .B(n242), .S(n505), .Z(n244) );
  MUX2_X1 U1435 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n511), .Z(n245) );
  MUX2_X1 U1436 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n510), .Z(n246) );
  MUX2_X1 U1437 ( .A(n246), .B(n245), .S(N11), .Z(n247) );
  MUX2_X1 U1438 ( .A(n247), .B(n244), .S(n500), .Z(n248) );
  MUX2_X1 U1439 ( .A(n248), .B(n241), .S(N13), .Z(n249) );
  MUX2_X1 U1440 ( .A(n249), .B(n234), .S(N14), .Z(n250) );
  MUX2_X1 U1441 ( .A(\mem[62][4] ), .B(\mem[63][4] ), .S(N10), .Z(n251) );
  MUX2_X1 U1442 ( .A(\mem[60][4] ), .B(\mem[61][4] ), .S(n512), .Z(n252) );
  MUX2_X1 U1443 ( .A(n252), .B(n251), .S(n503), .Z(n253) );
  MUX2_X1 U1444 ( .A(\mem[58][4] ), .B(\mem[59][4] ), .S(n512), .Z(n254) );
  MUX2_X1 U1445 ( .A(\mem[56][4] ), .B(\mem[57][4] ), .S(n512), .Z(n255) );
  MUX2_X1 U1446 ( .A(n255), .B(n254), .S(n503), .Z(n256) );
  MUX2_X1 U1447 ( .A(n256), .B(n253), .S(n500), .Z(n257) );
  MUX2_X1 U1448 ( .A(\mem[54][4] ), .B(\mem[55][4] ), .S(n512), .Z(n258) );
  MUX2_X1 U1449 ( .A(\mem[52][4] ), .B(\mem[53][4] ), .S(n513), .Z(n259) );
  MUX2_X1 U1450 ( .A(n259), .B(n258), .S(n504), .Z(n260) );
  MUX2_X1 U1451 ( .A(\mem[50][4] ), .B(\mem[51][4] ), .S(n512), .Z(n261) );
  MUX2_X1 U1452 ( .A(\mem[48][4] ), .B(\mem[49][4] ), .S(n512), .Z(n262) );
  MUX2_X1 U1453 ( .A(n262), .B(n261), .S(n504), .Z(n263) );
  MUX2_X1 U1454 ( .A(n263), .B(n260), .S(n500), .Z(n264) );
  MUX2_X1 U1455 ( .A(n264), .B(n257), .S(n499), .Z(n265) );
  MUX2_X1 U1456 ( .A(\mem[46][4] ), .B(\mem[47][4] ), .S(n512), .Z(n266) );
  MUX2_X1 U1457 ( .A(\mem[44][4] ), .B(\mem[45][4] ), .S(n513), .Z(n267) );
  MUX2_X1 U1458 ( .A(n267), .B(n266), .S(n504), .Z(n268) );
  MUX2_X1 U1459 ( .A(\mem[42][4] ), .B(\mem[43][4] ), .S(n511), .Z(n269) );
  MUX2_X1 U1460 ( .A(\mem[40][4] ), .B(\mem[41][4] ), .S(n510), .Z(n270) );
  MUX2_X1 U1461 ( .A(n270), .B(n269), .S(n503), .Z(n271) );
  MUX2_X1 U1462 ( .A(n271), .B(n268), .S(n500), .Z(n272) );
  MUX2_X1 U1463 ( .A(\mem[38][4] ), .B(\mem[39][4] ), .S(n511), .Z(n273) );
  MUX2_X1 U1464 ( .A(\mem[36][4] ), .B(\mem[37][4] ), .S(n510), .Z(n274) );
  MUX2_X1 U1465 ( .A(n274), .B(n273), .S(n504), .Z(n275) );
  MUX2_X1 U1466 ( .A(\mem[34][4] ), .B(\mem[35][4] ), .S(n511), .Z(n276) );
  MUX2_X1 U1467 ( .A(\mem[32][4] ), .B(\mem[33][4] ), .S(n512), .Z(n277) );
  MUX2_X1 U1468 ( .A(n277), .B(n276), .S(n504), .Z(n278) );
  MUX2_X1 U1469 ( .A(n278), .B(n275), .S(n500), .Z(n279) );
  MUX2_X1 U1470 ( .A(n279), .B(n272), .S(N13), .Z(n280) );
  MUX2_X1 U1471 ( .A(n280), .B(n265), .S(N14), .Z(n281) );
  MUX2_X1 U1472 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n512), .Z(n282) );
  MUX2_X1 U1473 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n511), .Z(n283) );
  MUX2_X1 U1474 ( .A(n283), .B(n282), .S(n503), .Z(n284) );
  MUX2_X1 U1475 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n511), .Z(n285) );
  MUX2_X1 U1476 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n512), .Z(n286) );
  MUX2_X1 U1477 ( .A(n286), .B(n285), .S(n504), .Z(n287) );
  MUX2_X1 U1478 ( .A(n287), .B(n284), .S(n500), .Z(n288) );
  MUX2_X1 U1479 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n510), .Z(n289) );
  MUX2_X1 U1480 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n513), .Z(n290) );
  MUX2_X1 U1481 ( .A(n290), .B(n289), .S(n503), .Z(n291) );
  MUX2_X1 U1482 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n513), .Z(n292) );
  MUX2_X1 U1483 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n510), .Z(n293) );
  MUX2_X1 U1484 ( .A(n293), .B(n292), .S(n503), .Z(n294) );
  MUX2_X1 U1485 ( .A(n294), .B(n291), .S(n500), .Z(n295) );
  MUX2_X1 U1486 ( .A(n295), .B(n288), .S(N13), .Z(n296) );
  MUX2_X1 U1487 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n510), .Z(n297) );
  MUX2_X1 U1488 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n511), .Z(n298) );
  MUX2_X1 U1489 ( .A(n298), .B(n297), .S(n503), .Z(n299) );
  MUX2_X1 U1490 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n511), .Z(n300) );
  MUX2_X1 U1491 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n511), .Z(n301) );
  MUX2_X1 U1492 ( .A(n301), .B(n300), .S(n503), .Z(n302) );
  MUX2_X1 U1493 ( .A(n302), .B(n299), .S(n500), .Z(n303) );
  MUX2_X1 U1494 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n512), .Z(n304) );
  MUX2_X1 U1495 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n512), .Z(n305) );
  MUX2_X1 U1496 ( .A(n305), .B(n304), .S(n504), .Z(n306) );
  MUX2_X1 U1497 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n510), .Z(n307) );
  MUX2_X1 U1498 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n510), .Z(n308) );
  MUX2_X1 U1499 ( .A(n308), .B(n307), .S(n504), .Z(n309) );
  MUX2_X1 U1500 ( .A(n309), .B(n306), .S(n500), .Z(n310) );
  MUX2_X1 U1501 ( .A(n310), .B(n303), .S(N13), .Z(n311) );
  MUX2_X1 U1502 ( .A(n311), .B(n296), .S(N14), .Z(n312) );
  MUX2_X1 U1503 ( .A(n312), .B(n281), .S(N15), .Z(N19) );
  MUX2_X1 U1504 ( .A(\mem[62][5] ), .B(\mem[63][5] ), .S(n513), .Z(n313) );
  MUX2_X1 U1505 ( .A(\mem[60][5] ), .B(\mem[61][5] ), .S(n513), .Z(n314) );
  MUX2_X1 U1506 ( .A(n314), .B(n313), .S(N11), .Z(n315) );
  MUX2_X1 U1507 ( .A(\mem[58][5] ), .B(\mem[59][5] ), .S(n513), .Z(n316) );
  MUX2_X1 U1508 ( .A(\mem[56][5] ), .B(\mem[57][5] ), .S(n513), .Z(n317) );
  MUX2_X1 U1509 ( .A(n317), .B(n316), .S(N11), .Z(n318) );
  MUX2_X1 U1510 ( .A(n318), .B(n315), .S(n501), .Z(n319) );
  MUX2_X1 U1511 ( .A(\mem[54][5] ), .B(\mem[55][5] ), .S(n513), .Z(n320) );
  MUX2_X1 U1512 ( .A(\mem[52][5] ), .B(\mem[53][5] ), .S(n513), .Z(n321) );
  MUX2_X1 U1513 ( .A(n321), .B(n320), .S(N11), .Z(n322) );
  MUX2_X1 U1514 ( .A(\mem[50][5] ), .B(\mem[51][5] ), .S(n513), .Z(n323) );
  MUX2_X1 U1515 ( .A(\mem[48][5] ), .B(\mem[49][5] ), .S(n512), .Z(n324) );
  MUX2_X1 U1516 ( .A(n324), .B(n323), .S(n509), .Z(n325) );
  MUX2_X1 U1517 ( .A(n325), .B(n322), .S(n501), .Z(n326) );
  MUX2_X1 U1518 ( .A(n326), .B(n319), .S(n499), .Z(n327) );
  MUX2_X1 U1519 ( .A(\mem[46][5] ), .B(\mem[47][5] ), .S(n513), .Z(n328) );
  MUX2_X1 U1520 ( .A(\mem[44][5] ), .B(\mem[45][5] ), .S(n513), .Z(n329) );
  MUX2_X1 U1521 ( .A(n329), .B(n328), .S(N11), .Z(n330) );
  MUX2_X1 U1522 ( .A(\mem[42][5] ), .B(\mem[43][5] ), .S(n513), .Z(n331) );
  MUX2_X1 U1523 ( .A(\mem[40][5] ), .B(\mem[41][5] ), .S(n511), .Z(n332) );
  MUX2_X1 U1524 ( .A(n332), .B(n331), .S(n509), .Z(n333) );
  MUX2_X1 U1525 ( .A(n333), .B(n330), .S(n501), .Z(n334) );
  MUX2_X1 U1526 ( .A(\mem[38][5] ), .B(\mem[39][5] ), .S(n516), .Z(n335) );
  MUX2_X1 U1527 ( .A(\mem[36][5] ), .B(\mem[37][5] ), .S(n512), .Z(n336) );
  MUX2_X1 U1528 ( .A(n336), .B(n335), .S(n509), .Z(n337) );
  MUX2_X1 U1529 ( .A(\mem[34][5] ), .B(\mem[35][5] ), .S(n510), .Z(n338) );
  MUX2_X1 U1530 ( .A(\mem[32][5] ), .B(\mem[33][5] ), .S(n512), .Z(n339) );
  MUX2_X1 U1531 ( .A(n339), .B(n338), .S(n509), .Z(n340) );
  MUX2_X1 U1532 ( .A(n340), .B(n337), .S(n501), .Z(n341) );
  MUX2_X1 U1533 ( .A(n341), .B(n334), .S(N13), .Z(n342) );
  MUX2_X1 U1534 ( .A(n342), .B(n327), .S(N14), .Z(n343) );
  MUX2_X1 U1535 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n510), .Z(n344) );
  MUX2_X1 U1536 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n510), .Z(n345) );
  MUX2_X1 U1537 ( .A(n345), .B(n344), .S(n507), .Z(n346) );
  MUX2_X1 U1538 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n513), .Z(n347) );
  MUX2_X1 U1539 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n512), .Z(n348) );
  MUX2_X1 U1540 ( .A(n348), .B(n347), .S(n509), .Z(n349) );
  MUX2_X1 U1541 ( .A(n349), .B(n346), .S(n501), .Z(n350) );
  MUX2_X1 U1542 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n512), .Z(n351) );
  MUX2_X1 U1543 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n512), .Z(n352) );
  MUX2_X1 U1544 ( .A(n352), .B(n351), .S(n506), .Z(n353) );
  MUX2_X1 U1545 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n511), .Z(n354) );
  MUX2_X1 U1546 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n511), .Z(n355) );
  MUX2_X1 U1547 ( .A(n355), .B(n354), .S(n509), .Z(n356) );
  MUX2_X1 U1548 ( .A(n356), .B(n353), .S(n501), .Z(n357) );
  MUX2_X1 U1549 ( .A(n357), .B(n350), .S(n499), .Z(n358) );
  MUX2_X1 U1550 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n510), .Z(n359) );
  MUX2_X1 U1551 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n511), .Z(n360) );
  MUX2_X1 U1552 ( .A(n360), .B(n359), .S(n506), .Z(n361) );
  MUX2_X1 U1553 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n515), .Z(n362) );
  MUX2_X1 U1554 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n510), .Z(n363) );
  MUX2_X1 U1555 ( .A(n363), .B(n362), .S(n506), .Z(n364) );
  MUX2_X1 U1556 ( .A(n364), .B(n361), .S(n501), .Z(n365) );
  MUX2_X1 U1557 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n1), .Z(n366) );
  MUX2_X1 U1558 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n513), .Z(n367) );
  MUX2_X1 U1559 ( .A(n367), .B(n366), .S(n506), .Z(n368) );
  MUX2_X1 U1560 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n515), .Z(n369) );
  MUX2_X1 U1561 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n511), .Z(n370) );
  MUX2_X1 U1562 ( .A(n370), .B(n369), .S(n506), .Z(n371) );
  MUX2_X1 U1563 ( .A(n371), .B(n368), .S(n501), .Z(n372) );
  MUX2_X1 U1564 ( .A(n372), .B(n365), .S(n499), .Z(n373) );
  MUX2_X1 U1565 ( .A(n373), .B(n358), .S(N14), .Z(n374) );
  MUX2_X1 U1566 ( .A(\mem[62][6] ), .B(\mem[63][6] ), .S(n511), .Z(n375) );
  MUX2_X1 U1567 ( .A(\mem[60][6] ), .B(\mem[61][6] ), .S(n511), .Z(n376) );
  MUX2_X1 U1568 ( .A(n376), .B(n375), .S(n506), .Z(n377) );
  MUX2_X1 U1569 ( .A(\mem[58][6] ), .B(\mem[59][6] ), .S(n514), .Z(n378) );
  MUX2_X1 U1570 ( .A(\mem[56][6] ), .B(\mem[57][6] ), .S(n515), .Z(n379) );
  MUX2_X1 U1571 ( .A(n379), .B(n378), .S(n506), .Z(n380) );
  MUX2_X1 U1572 ( .A(n380), .B(n377), .S(n501), .Z(n381) );
  MUX2_X1 U1573 ( .A(\mem[54][6] ), .B(\mem[55][6] ), .S(n1), .Z(n382) );
  MUX2_X1 U1574 ( .A(\mem[52][6] ), .B(\mem[53][6] ), .S(n512), .Z(n383) );
  MUX2_X1 U1575 ( .A(n383), .B(n382), .S(n506), .Z(n384) );
  MUX2_X1 U1576 ( .A(\mem[50][6] ), .B(\mem[51][6] ), .S(n1), .Z(n385) );
  MUX2_X1 U1577 ( .A(\mem[48][6] ), .B(\mem[49][6] ), .S(n1), .Z(n386) );
  MUX2_X1 U1578 ( .A(n386), .B(n385), .S(n506), .Z(n387) );
  MUX2_X1 U1579 ( .A(n387), .B(n384), .S(n501), .Z(n388) );
  MUX2_X1 U1580 ( .A(n388), .B(n381), .S(N13), .Z(n389) );
  MUX2_X1 U1581 ( .A(\mem[46][6] ), .B(\mem[47][6] ), .S(n511), .Z(n390) );
  MUX2_X1 U1582 ( .A(\mem[44][6] ), .B(\mem[45][6] ), .S(n514), .Z(n391) );
  MUX2_X1 U1583 ( .A(n391), .B(n390), .S(n506), .Z(n392) );
  MUX2_X1 U1584 ( .A(\mem[42][6] ), .B(\mem[43][6] ), .S(n510), .Z(n393) );
  MUX2_X1 U1585 ( .A(\mem[40][6] ), .B(\mem[41][6] ), .S(n515), .Z(n394) );
  MUX2_X1 U1586 ( .A(n394), .B(n393), .S(n506), .Z(n395) );
  MUX2_X1 U1587 ( .A(n395), .B(n392), .S(n501), .Z(n396) );
  MUX2_X1 U1588 ( .A(\mem[38][6] ), .B(\mem[39][6] ), .S(n514), .Z(n397) );
  MUX2_X1 U1589 ( .A(\mem[36][6] ), .B(\mem[37][6] ), .S(n514), .Z(n398) );
  MUX2_X1 U1590 ( .A(n398), .B(n397), .S(n506), .Z(n399) );
  MUX2_X1 U1591 ( .A(\mem[34][6] ), .B(\mem[35][6] ), .S(n511), .Z(n400) );
  MUX2_X1 U1592 ( .A(\mem[32][6] ), .B(\mem[33][6] ), .S(n512), .Z(n401) );
  MUX2_X1 U1593 ( .A(n401), .B(n400), .S(n506), .Z(n402) );
  MUX2_X1 U1594 ( .A(n402), .B(n399), .S(n501), .Z(n403) );
  MUX2_X1 U1595 ( .A(n403), .B(n396), .S(n499), .Z(n404) );
  MUX2_X1 U1596 ( .A(n404), .B(n389), .S(N14), .Z(n405) );
  MUX2_X1 U1597 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n515), .Z(n406) );
  MUX2_X1 U1598 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n515), .Z(n407) );
  MUX2_X1 U1599 ( .A(n407), .B(n406), .S(n507), .Z(n408) );
  MUX2_X1 U1600 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n516), .Z(n409) );
  MUX2_X1 U1601 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n510), .Z(n410) );
  MUX2_X1 U1602 ( .A(n410), .B(n409), .S(n507), .Z(n411) );
  MUX2_X1 U1603 ( .A(n411), .B(n408), .S(n502), .Z(n412) );
  MUX2_X1 U1604 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n516), .Z(n413) );
  MUX2_X1 U1605 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n515), .Z(n414) );
  MUX2_X1 U1606 ( .A(n414), .B(n413), .S(n507), .Z(n415) );
  MUX2_X1 U1607 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n513), .Z(n416) );
  MUX2_X1 U1608 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n515), .Z(n417) );
  MUX2_X1 U1609 ( .A(n417), .B(n416), .S(n507), .Z(n418) );
  MUX2_X1 U1610 ( .A(n418), .B(n415), .S(n502), .Z(n419) );
  MUX2_X1 U1611 ( .A(n419), .B(n412), .S(n499), .Z(n420) );
  MUX2_X1 U1612 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n514), .Z(n421) );
  MUX2_X1 U1613 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n514), .Z(n422) );
  MUX2_X1 U1614 ( .A(n422), .B(n421), .S(n507), .Z(n423) );
  MUX2_X1 U1615 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n516), .Z(n424) );
  MUX2_X1 U1616 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n514), .Z(n425) );
  MUX2_X1 U1617 ( .A(n425), .B(n424), .S(n507), .Z(n426) );
  MUX2_X1 U1618 ( .A(n426), .B(n423), .S(n502), .Z(n427) );
  MUX2_X1 U1619 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n513), .Z(n428) );
  MUX2_X1 U1620 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n512), .Z(n429) );
  MUX2_X1 U1621 ( .A(n429), .B(n428), .S(n507), .Z(n430) );
  MUX2_X1 U1622 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n511), .Z(n431) );
  MUX2_X1 U1623 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n1), .Z(n432) );
  MUX2_X1 U1624 ( .A(n432), .B(n431), .S(n507), .Z(n433) );
  MUX2_X1 U1625 ( .A(n433), .B(n430), .S(n502), .Z(n434) );
  MUX2_X1 U1626 ( .A(n434), .B(n427), .S(n499), .Z(n435) );
  MUX2_X1 U1627 ( .A(n435), .B(n420), .S(N14), .Z(n436) );
  MUX2_X1 U1628 ( .A(\mem[62][7] ), .B(\mem[63][7] ), .S(n516), .Z(n437) );
  MUX2_X1 U1629 ( .A(\mem[60][7] ), .B(\mem[61][7] ), .S(n510), .Z(n438) );
  MUX2_X1 U1630 ( .A(n438), .B(n437), .S(n507), .Z(n439) );
  MUX2_X1 U1631 ( .A(\mem[58][7] ), .B(\mem[59][7] ), .S(n514), .Z(n440) );
  MUX2_X1 U1632 ( .A(\mem[56][7] ), .B(\mem[57][7] ), .S(n1), .Z(n441) );
  MUX2_X1 U1633 ( .A(n441), .B(n440), .S(n507), .Z(n442) );
  MUX2_X1 U1634 ( .A(n442), .B(n439), .S(n502), .Z(n443) );
  MUX2_X1 U1635 ( .A(\mem[54][7] ), .B(\mem[55][7] ), .S(n1), .Z(n444) );
  MUX2_X1 U1636 ( .A(\mem[52][7] ), .B(\mem[53][7] ), .S(n512), .Z(n445) );
  MUX2_X1 U1637 ( .A(n445), .B(n444), .S(n507), .Z(n446) );
  MUX2_X1 U1638 ( .A(\mem[50][7] ), .B(\mem[51][7] ), .S(n515), .Z(n447) );
  MUX2_X1 U1639 ( .A(\mem[48][7] ), .B(\mem[49][7] ), .S(n515), .Z(n448) );
  MUX2_X1 U1640 ( .A(n448), .B(n447), .S(n507), .Z(n449) );
  MUX2_X1 U1641 ( .A(n449), .B(n446), .S(n502), .Z(n450) );
  MUX2_X1 U1642 ( .A(n450), .B(n443), .S(n499), .Z(n451) );
  MUX2_X1 U1643 ( .A(\mem[46][7] ), .B(\mem[47][7] ), .S(n510), .Z(n452) );
  MUX2_X1 U1644 ( .A(\mem[44][7] ), .B(\mem[45][7] ), .S(n511), .Z(n453) );
  MUX2_X1 U1645 ( .A(n453), .B(n452), .S(n508), .Z(n454) );
  MUX2_X1 U1646 ( .A(\mem[42][7] ), .B(\mem[43][7] ), .S(n511), .Z(n455) );
  MUX2_X1 U1647 ( .A(\mem[40][7] ), .B(\mem[41][7] ), .S(n511), .Z(n456) );
  MUX2_X1 U1648 ( .A(n456), .B(n455), .S(n508), .Z(n457) );
  MUX2_X1 U1649 ( .A(n457), .B(n454), .S(n502), .Z(n458) );
  MUX2_X1 U1650 ( .A(\mem[38][7] ), .B(\mem[39][7] ), .S(n516), .Z(n459) );
  MUX2_X1 U1651 ( .A(\mem[36][7] ), .B(\mem[37][7] ), .S(n513), .Z(n460) );
  MUX2_X1 U1652 ( .A(n460), .B(n459), .S(n508), .Z(n461) );
  MUX2_X1 U1653 ( .A(\mem[34][7] ), .B(\mem[35][7] ), .S(n513), .Z(n462) );
  MUX2_X1 U1654 ( .A(\mem[32][7] ), .B(\mem[33][7] ), .S(n510), .Z(n463) );
  MUX2_X1 U1655 ( .A(n463), .B(n462), .S(n508), .Z(n464) );
  MUX2_X1 U1656 ( .A(n464), .B(n461), .S(n502), .Z(n465) );
  MUX2_X1 U1657 ( .A(n465), .B(n458), .S(N13), .Z(n466) );
  MUX2_X1 U1658 ( .A(n466), .B(n451), .S(N14), .Z(n467) );
  MUX2_X1 U1659 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n511), .Z(n468) );
  MUX2_X1 U1660 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n513), .Z(n469) );
  MUX2_X1 U1661 ( .A(n469), .B(n468), .S(n508), .Z(n470) );
  MUX2_X1 U1662 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n516), .Z(n471) );
  MUX2_X1 U1663 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n510), .Z(n472) );
  MUX2_X1 U1664 ( .A(n472), .B(n471), .S(n508), .Z(n473) );
  MUX2_X1 U1665 ( .A(n473), .B(n470), .S(n502), .Z(n474) );
  MUX2_X1 U1666 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n512), .Z(n475) );
  MUX2_X1 U1667 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n511), .Z(n476) );
  MUX2_X1 U1668 ( .A(n476), .B(n475), .S(n508), .Z(n477) );
  MUX2_X1 U1669 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n1), .Z(n478) );
  MUX2_X1 U1670 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n512), .Z(n479) );
  MUX2_X1 U1671 ( .A(n479), .B(n478), .S(n508), .Z(n480) );
  MUX2_X1 U1672 ( .A(n480), .B(n477), .S(n502), .Z(n481) );
  MUX2_X1 U1673 ( .A(n481), .B(n474), .S(n499), .Z(n482) );
  MUX2_X1 U1674 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n1), .Z(n483) );
  MUX2_X1 U1675 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n1), .Z(n484) );
  MUX2_X1 U1676 ( .A(n484), .B(n483), .S(n508), .Z(n485) );
  MUX2_X1 U1677 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n512), .Z(n486) );
  MUX2_X1 U1678 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n511), .Z(n487) );
  MUX2_X1 U1679 ( .A(n487), .B(n486), .S(n508), .Z(n488) );
  MUX2_X1 U1680 ( .A(n488), .B(n485), .S(n502), .Z(n489) );
  MUX2_X1 U1681 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n514), .Z(n490) );
  MUX2_X1 U1682 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n1), .Z(n491) );
  MUX2_X1 U1683 ( .A(n491), .B(n490), .S(n508), .Z(n492) );
  MUX2_X1 U1684 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n514), .Z(n493) );
  MUX2_X1 U1685 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n515), .Z(n494) );
  MUX2_X1 U1686 ( .A(n494), .B(n493), .S(n508), .Z(n495) );
  MUX2_X1 U1687 ( .A(n495), .B(n492), .S(n502), .Z(n496) );
  MUX2_X1 U1688 ( .A(n496), .B(n489), .S(N13), .Z(n497) );
  MUX2_X1 U1689 ( .A(n497), .B(n482), .S(N14), .Z(n498) );
  CLKBUF_X1 U1690 ( .A(N12), .Z(n500) );
  CLKBUF_X1 U1691 ( .A(N12), .Z(n502) );
  INV_X1 U1692 ( .A(N10), .ZN(n518) );
  INV_X1 U1693 ( .A(N11), .ZN(n519) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N15), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N17), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N19), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N21), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N23), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N25), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N27), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n285), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n284), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n283), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n282), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n281), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n280), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n279), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n278), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n277), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n276), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n275), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n274), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n273), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n272), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n271), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n270), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n269), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n268), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n267), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n266), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n265), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n264), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n263), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n262), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n261), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n260), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n259), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n258), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n257), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n256), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n255), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n254), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n253), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n252), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n251), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n250), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n249), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n248), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n247), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n246), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n245), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n244), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n243), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n242), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n241), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n240), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n239), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n238), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n237), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n236), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n235), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n234), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n233), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n232), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n231), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n230), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n229), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n228), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n227), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n226), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n225), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n224), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n223), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n222), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n221), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n220), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n219), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n218), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n217), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n216), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n215), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n214), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n213), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n212), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n211), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n210), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n209), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n208), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n207), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n206), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n205), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n204), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n203), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n202), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n201), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n200), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n199), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n198), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n197), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n196), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n195), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n194), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n193), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n192), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n191), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n190), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n189), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n188), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n187), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n186), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n185), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n184), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n183), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n182), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n181), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n180), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n179), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n178), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n177), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n176), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n175), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n174), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n173), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n172), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n171), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n170), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n169), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n168), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n167), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n166), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n165), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n164), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n163), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n162), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n161), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n160), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n159), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n158), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n37), .ZN(n20) );
  NAND3_X1 U281 ( .A1(n37), .A2(n376), .A3(N10), .ZN(n38) );
  NAND3_X1 U282 ( .A1(n37), .A2(n375), .A3(N11), .ZN(n55) );
  NAND3_X1 U283 ( .A1(N10), .A2(n37), .A3(N11), .ZN(n72) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n106), .ZN(n89) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n106), .ZN(n107) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n106), .ZN(n124) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n106), .ZN(n141) );
  BUF_X1 U3 ( .A(N10), .Z(n365) );
  BUF_X1 U4 ( .A(N10), .Z(n366) );
  BUF_X1 U5 ( .A(n20), .Z(n374) );
  BUF_X1 U6 ( .A(n38), .Z(n373) );
  BUF_X1 U7 ( .A(n55), .Z(n372) );
  BUF_X1 U8 ( .A(n72), .Z(n371) );
  BUF_X1 U9 ( .A(n124), .Z(n368) );
  BUF_X1 U10 ( .A(n141), .Z(n367) );
  BUF_X1 U11 ( .A(n89), .Z(n370) );
  BUF_X1 U12 ( .A(n107), .Z(n369) );
  BUF_X1 U13 ( .A(N10), .Z(n364) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  INV_X1 U15 ( .A(data_in[4]), .ZN(n382) );
  INV_X1 U16 ( .A(data_in[5]), .ZN(n383) );
  INV_X1 U17 ( .A(data_in[6]), .ZN(n384) );
  INV_X1 U18 ( .A(data_in[7]), .ZN(n385) );
  INV_X1 U19 ( .A(data_in[8]), .ZN(n386) );
  INV_X1 U20 ( .A(data_in[9]), .ZN(n387) );
  INV_X1 U21 ( .A(data_in[11]), .ZN(n389) );
  INV_X1 U22 ( .A(data_in[12]), .ZN(n390) );
  INV_X1 U23 ( .A(data_in[13]), .ZN(n391) );
  INV_X1 U24 ( .A(data_in[1]), .ZN(n379) );
  INV_X1 U25 ( .A(data_in[2]), .ZN(n380) );
  INV_X1 U26 ( .A(data_in[3]), .ZN(n381) );
  INV_X1 U27 ( .A(data_in[10]), .ZN(n388) );
  INV_X1 U28 ( .A(data_in[14]), .ZN(n392) );
  INV_X1 U29 ( .A(data_in[15]), .ZN(n393) );
  NOR2_X1 U30 ( .A1(n377), .A2(N12), .ZN(n37) );
  INV_X1 U31 ( .A(wr_en), .ZN(n377) );
  OAI21_X1 U32 ( .B1(n374), .B2(n378), .A(n21), .ZN(n158) );
  NAND2_X1 U33 ( .A1(\mem[0][0] ), .A2(n20), .ZN(n21) );
  OAI21_X1 U34 ( .B1(n378), .B2(n38), .A(n39), .ZN(n174) );
  NAND2_X1 U35 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n39) );
  OAI21_X1 U36 ( .B1(n378), .B2(n55), .A(n56), .ZN(n190) );
  NAND2_X1 U37 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n56) );
  OAI21_X1 U38 ( .B1(n378), .B2(n72), .A(n73), .ZN(n206) );
  NAND2_X1 U39 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n73) );
  OAI21_X1 U40 ( .B1(n378), .B2(n370), .A(n90), .ZN(n222) );
  NAND2_X1 U41 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n90) );
  OAI21_X1 U42 ( .B1(n378), .B2(n369), .A(n108), .ZN(n238) );
  NAND2_X1 U43 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n108) );
  OAI21_X1 U44 ( .B1(n378), .B2(n124), .A(n125), .ZN(n254) );
  NAND2_X1 U45 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n125) );
  OAI21_X1 U46 ( .B1(n378), .B2(n141), .A(n142), .ZN(n270) );
  NAND2_X1 U47 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n142) );
  AND2_X1 U48 ( .A1(N12), .A2(wr_en), .ZN(n106) );
  INV_X1 U49 ( .A(N10), .ZN(n375) );
  OAI21_X1 U50 ( .B1(n385), .B2(n72), .A(n80), .ZN(n213) );
  NAND2_X1 U51 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n80) );
  OAI21_X1 U52 ( .B1(n386), .B2(n371), .A(n81), .ZN(n214) );
  NAND2_X1 U53 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n81) );
  OAI21_X1 U54 ( .B1(n387), .B2(n72), .A(n82), .ZN(n215) );
  NAND2_X1 U55 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n82) );
  OAI21_X1 U56 ( .B1(n388), .B2(n72), .A(n83), .ZN(n216) );
  NAND2_X1 U57 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n83) );
  OAI21_X1 U58 ( .B1(n389), .B2(n72), .A(n84), .ZN(n217) );
  NAND2_X1 U59 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n84) );
  OAI21_X1 U60 ( .B1(n390), .B2(n72), .A(n85), .ZN(n218) );
  NAND2_X1 U61 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n85) );
  OAI21_X1 U62 ( .B1(n391), .B2(n72), .A(n86), .ZN(n219) );
  NAND2_X1 U63 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n86) );
  OAI21_X1 U64 ( .B1(n392), .B2(n72), .A(n87), .ZN(n220) );
  NAND2_X1 U65 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n87) );
  OAI21_X1 U66 ( .B1(n385), .B2(n107), .A(n115), .ZN(n245) );
  NAND2_X1 U67 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n115) );
  OAI21_X1 U68 ( .B1(n386), .B2(n107), .A(n116), .ZN(n246) );
  NAND2_X1 U69 ( .A1(\mem[5][8] ), .A2(n107), .ZN(n116) );
  OAI21_X1 U70 ( .B1(n387), .B2(n107), .A(n117), .ZN(n247) );
  NAND2_X1 U71 ( .A1(\mem[5][9] ), .A2(n107), .ZN(n117) );
  OAI21_X1 U72 ( .B1(n388), .B2(n107), .A(n118), .ZN(n248) );
  NAND2_X1 U73 ( .A1(\mem[5][10] ), .A2(n107), .ZN(n118) );
  OAI21_X1 U74 ( .B1(n389), .B2(n107), .A(n119), .ZN(n249) );
  NAND2_X1 U75 ( .A1(\mem[5][11] ), .A2(n107), .ZN(n119) );
  OAI21_X1 U76 ( .B1(n390), .B2(n107), .A(n120), .ZN(n250) );
  NAND2_X1 U77 ( .A1(\mem[5][12] ), .A2(n107), .ZN(n120) );
  OAI21_X1 U78 ( .B1(n391), .B2(n107), .A(n121), .ZN(n251) );
  NAND2_X1 U79 ( .A1(\mem[5][13] ), .A2(n107), .ZN(n121) );
  OAI21_X1 U80 ( .B1(n392), .B2(n107), .A(n122), .ZN(n252) );
  NAND2_X1 U81 ( .A1(\mem[5][14] ), .A2(n107), .ZN(n122) );
  OAI21_X1 U82 ( .B1(n385), .B2(n141), .A(n149), .ZN(n277) );
  NAND2_X1 U83 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n149) );
  OAI21_X1 U84 ( .B1(n386), .B2(n141), .A(n150), .ZN(n278) );
  NAND2_X1 U85 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n150) );
  OAI21_X1 U86 ( .B1(n387), .B2(n367), .A(n151), .ZN(n279) );
  NAND2_X1 U87 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n151) );
  OAI21_X1 U88 ( .B1(n388), .B2(n141), .A(n152), .ZN(n280) );
  NAND2_X1 U89 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n152) );
  OAI21_X1 U90 ( .B1(n389), .B2(n141), .A(n153), .ZN(n281) );
  NAND2_X1 U91 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n153) );
  OAI21_X1 U92 ( .B1(n390), .B2(n141), .A(n154), .ZN(n282) );
  NAND2_X1 U93 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n154) );
  OAI21_X1 U94 ( .B1(n391), .B2(n141), .A(n155), .ZN(n283) );
  NAND2_X1 U95 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n155) );
  OAI21_X1 U96 ( .B1(n392), .B2(n141), .A(n156), .ZN(n284) );
  NAND2_X1 U97 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n156) );
  OAI21_X1 U98 ( .B1(n385), .B2(n38), .A(n46), .ZN(n181) );
  NAND2_X1 U99 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n46) );
  OAI21_X1 U100 ( .B1(n386), .B2(n373), .A(n47), .ZN(n182) );
  NAND2_X1 U101 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n47) );
  OAI21_X1 U102 ( .B1(n387), .B2(n38), .A(n48), .ZN(n183) );
  NAND2_X1 U103 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n48) );
  OAI21_X1 U104 ( .B1(n388), .B2(n38), .A(n49), .ZN(n184) );
  NAND2_X1 U105 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n49) );
  OAI21_X1 U106 ( .B1(n389), .B2(n38), .A(n50), .ZN(n185) );
  NAND2_X1 U107 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n50) );
  OAI21_X1 U108 ( .B1(n390), .B2(n38), .A(n51), .ZN(n186) );
  NAND2_X1 U109 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n51) );
  OAI21_X1 U110 ( .B1(n391), .B2(n38), .A(n52), .ZN(n187) );
  NAND2_X1 U111 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n52) );
  OAI21_X1 U112 ( .B1(n392), .B2(n38), .A(n53), .ZN(n188) );
  NAND2_X1 U113 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n53) );
  OAI21_X1 U114 ( .B1(n385), .B2(n124), .A(n132), .ZN(n261) );
  NAND2_X1 U115 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n132) );
  OAI21_X1 U116 ( .B1(n386), .B2(n368), .A(n133), .ZN(n262) );
  NAND2_X1 U117 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n133) );
  OAI21_X1 U118 ( .B1(n387), .B2(n124), .A(n134), .ZN(n263) );
  NAND2_X1 U119 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n134) );
  OAI21_X1 U120 ( .B1(n388), .B2(n124), .A(n135), .ZN(n264) );
  NAND2_X1 U121 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n135) );
  OAI21_X1 U122 ( .B1(n389), .B2(n124), .A(n136), .ZN(n265) );
  NAND2_X1 U123 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n136) );
  OAI21_X1 U124 ( .B1(n390), .B2(n124), .A(n137), .ZN(n266) );
  NAND2_X1 U125 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n137) );
  OAI21_X1 U126 ( .B1(n391), .B2(n124), .A(n138), .ZN(n267) );
  NAND2_X1 U127 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n138) );
  OAI21_X1 U128 ( .B1(n392), .B2(n124), .A(n139), .ZN(n268) );
  NAND2_X1 U129 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n139) );
  OAI21_X1 U130 ( .B1(n385), .B2(n55), .A(n63), .ZN(n197) );
  NAND2_X1 U131 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n63) );
  OAI21_X1 U132 ( .B1(n386), .B2(n372), .A(n64), .ZN(n198) );
  NAND2_X1 U133 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n64) );
  OAI21_X1 U134 ( .B1(n387), .B2(n55), .A(n65), .ZN(n199) );
  NAND2_X1 U135 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n65) );
  OAI21_X1 U136 ( .B1(n388), .B2(n55), .A(n66), .ZN(n200) );
  NAND2_X1 U137 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n66) );
  OAI21_X1 U138 ( .B1(n389), .B2(n55), .A(n67), .ZN(n201) );
  NAND2_X1 U139 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n67) );
  OAI21_X1 U140 ( .B1(n390), .B2(n55), .A(n68), .ZN(n202) );
  NAND2_X1 U141 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n68) );
  OAI21_X1 U142 ( .B1(n391), .B2(n55), .A(n69), .ZN(n203) );
  NAND2_X1 U143 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n69) );
  OAI21_X1 U144 ( .B1(n392), .B2(n55), .A(n70), .ZN(n204) );
  NAND2_X1 U145 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n70) );
  OAI21_X1 U146 ( .B1(n385), .B2(n89), .A(n97), .ZN(n229) );
  NAND2_X1 U147 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n97) );
  OAI21_X1 U148 ( .B1(n386), .B2(n89), .A(n98), .ZN(n230) );
  NAND2_X1 U149 ( .A1(\mem[4][8] ), .A2(n89), .ZN(n98) );
  OAI21_X1 U150 ( .B1(n387), .B2(n89), .A(n99), .ZN(n231) );
  NAND2_X1 U151 ( .A1(\mem[4][9] ), .A2(n89), .ZN(n99) );
  OAI21_X1 U152 ( .B1(n388), .B2(n89), .A(n100), .ZN(n232) );
  NAND2_X1 U153 ( .A1(\mem[4][10] ), .A2(n89), .ZN(n100) );
  OAI21_X1 U154 ( .B1(n389), .B2(n89), .A(n101), .ZN(n233) );
  NAND2_X1 U155 ( .A1(\mem[4][11] ), .A2(n89), .ZN(n101) );
  OAI21_X1 U156 ( .B1(n390), .B2(n89), .A(n102), .ZN(n234) );
  NAND2_X1 U157 ( .A1(\mem[4][12] ), .A2(n89), .ZN(n102) );
  OAI21_X1 U158 ( .B1(n391), .B2(n89), .A(n103), .ZN(n235) );
  NAND2_X1 U159 ( .A1(\mem[4][13] ), .A2(n89), .ZN(n103) );
  OAI21_X1 U160 ( .B1(n392), .B2(n89), .A(n104), .ZN(n236) );
  NAND2_X1 U161 ( .A1(\mem[4][14] ), .A2(n89), .ZN(n104) );
  OAI21_X1 U162 ( .B1(n382), .B2(n38), .A(n43), .ZN(n178) );
  NAND2_X1 U163 ( .A1(\mem[1][4] ), .A2(n38), .ZN(n43) );
  OAI21_X1 U164 ( .B1(n383), .B2(n38), .A(n44), .ZN(n179) );
  NAND2_X1 U165 ( .A1(\mem[1][5] ), .A2(n38), .ZN(n44) );
  OAI21_X1 U166 ( .B1(n384), .B2(n38), .A(n45), .ZN(n180) );
  NAND2_X1 U167 ( .A1(\mem[1][6] ), .A2(n38), .ZN(n45) );
  OAI21_X1 U168 ( .B1(n382), .B2(n55), .A(n60), .ZN(n194) );
  NAND2_X1 U169 ( .A1(\mem[2][4] ), .A2(n55), .ZN(n60) );
  OAI21_X1 U170 ( .B1(n383), .B2(n55), .A(n61), .ZN(n195) );
  NAND2_X1 U171 ( .A1(\mem[2][5] ), .A2(n55), .ZN(n61) );
  OAI21_X1 U172 ( .B1(n384), .B2(n55), .A(n62), .ZN(n196) );
  NAND2_X1 U173 ( .A1(\mem[2][6] ), .A2(n55), .ZN(n62) );
  OAI21_X1 U174 ( .B1(n382), .B2(n72), .A(n77), .ZN(n210) );
  NAND2_X1 U175 ( .A1(\mem[3][4] ), .A2(n72), .ZN(n77) );
  OAI21_X1 U176 ( .B1(n383), .B2(n72), .A(n78), .ZN(n211) );
  NAND2_X1 U177 ( .A1(\mem[3][5] ), .A2(n72), .ZN(n78) );
  OAI21_X1 U178 ( .B1(n384), .B2(n72), .A(n79), .ZN(n212) );
  NAND2_X1 U179 ( .A1(\mem[3][6] ), .A2(n72), .ZN(n79) );
  OAI21_X1 U180 ( .B1(n382), .B2(n370), .A(n94), .ZN(n226) );
  NAND2_X1 U181 ( .A1(\mem[4][4] ), .A2(n370), .ZN(n94) );
  OAI21_X1 U182 ( .B1(n383), .B2(n370), .A(n95), .ZN(n227) );
  NAND2_X1 U183 ( .A1(\mem[4][5] ), .A2(n370), .ZN(n95) );
  OAI21_X1 U184 ( .B1(n384), .B2(n370), .A(n96), .ZN(n228) );
  NAND2_X1 U185 ( .A1(\mem[4][6] ), .A2(n370), .ZN(n96) );
  OAI21_X1 U186 ( .B1(n382), .B2(n369), .A(n112), .ZN(n242) );
  NAND2_X1 U187 ( .A1(\mem[5][4] ), .A2(n369), .ZN(n112) );
  OAI21_X1 U188 ( .B1(n383), .B2(n369), .A(n113), .ZN(n243) );
  NAND2_X1 U189 ( .A1(\mem[5][5] ), .A2(n369), .ZN(n113) );
  OAI21_X1 U190 ( .B1(n384), .B2(n369), .A(n114), .ZN(n244) );
  NAND2_X1 U191 ( .A1(\mem[5][6] ), .A2(n369), .ZN(n114) );
  OAI21_X1 U192 ( .B1(n382), .B2(n124), .A(n129), .ZN(n258) );
  NAND2_X1 U193 ( .A1(\mem[6][4] ), .A2(n124), .ZN(n129) );
  OAI21_X1 U194 ( .B1(n383), .B2(n124), .A(n130), .ZN(n259) );
  NAND2_X1 U195 ( .A1(\mem[6][5] ), .A2(n124), .ZN(n130) );
  OAI21_X1 U196 ( .B1(n384), .B2(n124), .A(n131), .ZN(n260) );
  NAND2_X1 U197 ( .A1(\mem[6][6] ), .A2(n124), .ZN(n131) );
  OAI21_X1 U198 ( .B1(n382), .B2(n141), .A(n146), .ZN(n274) );
  NAND2_X1 U199 ( .A1(\mem[7][4] ), .A2(n141), .ZN(n146) );
  OAI21_X1 U200 ( .B1(n383), .B2(n141), .A(n147), .ZN(n275) );
  NAND2_X1 U201 ( .A1(\mem[7][5] ), .A2(n141), .ZN(n147) );
  OAI21_X1 U202 ( .B1(n384), .B2(n141), .A(n148), .ZN(n276) );
  NAND2_X1 U203 ( .A1(\mem[7][6] ), .A2(n141), .ZN(n148) );
  OAI21_X1 U204 ( .B1(n20), .B2(n386), .A(n29), .ZN(n166) );
  NAND2_X1 U205 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n29) );
  OAI21_X1 U206 ( .B1(n20), .B2(n387), .A(n30), .ZN(n167) );
  NAND2_X1 U207 ( .A1(\mem[0][9] ), .A2(n20), .ZN(n30) );
  OAI21_X1 U208 ( .B1(n20), .B2(n388), .A(n31), .ZN(n168) );
  NAND2_X1 U209 ( .A1(\mem[0][10] ), .A2(n20), .ZN(n31) );
  OAI21_X1 U210 ( .B1(n20), .B2(n389), .A(n32), .ZN(n169) );
  NAND2_X1 U211 ( .A1(\mem[0][11] ), .A2(n20), .ZN(n32) );
  OAI21_X1 U212 ( .B1(n374), .B2(n390), .A(n33), .ZN(n170) );
  NAND2_X1 U213 ( .A1(\mem[0][12] ), .A2(n20), .ZN(n33) );
  OAI21_X1 U214 ( .B1(n20), .B2(n391), .A(n34), .ZN(n171) );
  NAND2_X1 U215 ( .A1(\mem[0][13] ), .A2(n20), .ZN(n34) );
  OAI21_X1 U216 ( .B1(n20), .B2(n392), .A(n35), .ZN(n172) );
  NAND2_X1 U217 ( .A1(\mem[0][14] ), .A2(n20), .ZN(n35) );
  INV_X1 U218 ( .A(N11), .ZN(n376) );
  OAI21_X1 U219 ( .B1(n374), .B2(n382), .A(n25), .ZN(n162) );
  NAND2_X1 U220 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n25) );
  OAI21_X1 U221 ( .B1(n374), .B2(n383), .A(n26), .ZN(n163) );
  NAND2_X1 U222 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n26) );
  OAI21_X1 U223 ( .B1(n374), .B2(n384), .A(n27), .ZN(n164) );
  NAND2_X1 U224 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n27) );
  OAI21_X1 U225 ( .B1(n374), .B2(n385), .A(n28), .ZN(n165) );
  NAND2_X1 U226 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n28) );
  OAI21_X1 U227 ( .B1(n379), .B2(n38), .A(n40), .ZN(n175) );
  NAND2_X1 U228 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n40) );
  OAI21_X1 U229 ( .B1(n381), .B2(n38), .A(n42), .ZN(n177) );
  NAND2_X1 U230 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n42) );
  OAI21_X1 U231 ( .B1(n379), .B2(n55), .A(n57), .ZN(n191) );
  NAND2_X1 U232 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n57) );
  OAI21_X1 U233 ( .B1(n381), .B2(n55), .A(n59), .ZN(n193) );
  NAND2_X1 U234 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n59) );
  OAI21_X1 U235 ( .B1(n379), .B2(n72), .A(n74), .ZN(n207) );
  NAND2_X1 U236 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n74) );
  OAI21_X1 U237 ( .B1(n381), .B2(n72), .A(n76), .ZN(n209) );
  NAND2_X1 U238 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n76) );
  OAI21_X1 U239 ( .B1(n379), .B2(n370), .A(n91), .ZN(n223) );
  NAND2_X1 U240 ( .A1(\mem[4][1] ), .A2(n89), .ZN(n91) );
  OAI21_X1 U241 ( .B1(n381), .B2(n370), .A(n93), .ZN(n225) );
  NAND2_X1 U242 ( .A1(\mem[4][3] ), .A2(n89), .ZN(n93) );
  OAI21_X1 U243 ( .B1(n379), .B2(n369), .A(n109), .ZN(n239) );
  NAND2_X1 U244 ( .A1(\mem[5][1] ), .A2(n107), .ZN(n109) );
  OAI21_X1 U245 ( .B1(n381), .B2(n369), .A(n111), .ZN(n241) );
  NAND2_X1 U246 ( .A1(\mem[5][3] ), .A2(n107), .ZN(n111) );
  OAI21_X1 U247 ( .B1(n379), .B2(n124), .A(n126), .ZN(n255) );
  NAND2_X1 U248 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n126) );
  OAI21_X1 U249 ( .B1(n381), .B2(n124), .A(n128), .ZN(n257) );
  NAND2_X1 U250 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n128) );
  OAI21_X1 U251 ( .B1(n379), .B2(n141), .A(n143), .ZN(n271) );
  NAND2_X1 U252 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n143) );
  OAI21_X1 U253 ( .B1(n381), .B2(n141), .A(n145), .ZN(n273) );
  NAND2_X1 U254 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n145) );
  OAI21_X1 U255 ( .B1(n380), .B2(n38), .A(n41), .ZN(n176) );
  NAND2_X1 U256 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n41) );
  OAI21_X1 U257 ( .B1(n380), .B2(n55), .A(n58), .ZN(n192) );
  NAND2_X1 U258 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n58) );
  OAI21_X1 U259 ( .B1(n380), .B2(n72), .A(n75), .ZN(n208) );
  NAND2_X1 U260 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n75) );
  OAI21_X1 U261 ( .B1(n380), .B2(n370), .A(n92), .ZN(n224) );
  NAND2_X1 U262 ( .A1(\mem[4][2] ), .A2(n89), .ZN(n92) );
  OAI21_X1 U263 ( .B1(n380), .B2(n369), .A(n110), .ZN(n240) );
  NAND2_X1 U264 ( .A1(\mem[5][2] ), .A2(n107), .ZN(n110) );
  OAI21_X1 U265 ( .B1(n380), .B2(n124), .A(n127), .ZN(n256) );
  NAND2_X1 U266 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n127) );
  OAI21_X1 U267 ( .B1(n380), .B2(n141), .A(n144), .ZN(n272) );
  NAND2_X1 U268 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n144) );
  OAI21_X1 U269 ( .B1(n393), .B2(n38), .A(n54), .ZN(n189) );
  NAND2_X1 U270 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n54) );
  OAI21_X1 U271 ( .B1(n393), .B2(n55), .A(n71), .ZN(n205) );
  NAND2_X1 U272 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n71) );
  OAI21_X1 U273 ( .B1(n393), .B2(n72), .A(n88), .ZN(n221) );
  NAND2_X1 U274 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n88) );
  OAI21_X1 U275 ( .B1(n393), .B2(n370), .A(n105), .ZN(n237) );
  NAND2_X1 U276 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n105) );
  OAI21_X1 U277 ( .B1(n393), .B2(n369), .A(n123), .ZN(n253) );
  NAND2_X1 U278 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n123) );
  OAI21_X1 U279 ( .B1(n393), .B2(n124), .A(n140), .ZN(n269) );
  NAND2_X1 U288 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n140) );
  OAI21_X1 U289 ( .B1(n393), .B2(n141), .A(n157), .ZN(n285) );
  NAND2_X1 U290 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n157) );
  OAI21_X1 U291 ( .B1(n374), .B2(n379), .A(n22), .ZN(n159) );
  NAND2_X1 U292 ( .A1(\mem[0][1] ), .A2(n20), .ZN(n22) );
  OAI21_X1 U293 ( .B1(n374), .B2(n380), .A(n23), .ZN(n160) );
  NAND2_X1 U294 ( .A1(\mem[0][2] ), .A2(n20), .ZN(n23) );
  OAI21_X1 U295 ( .B1(n374), .B2(n381), .A(n24), .ZN(n161) );
  NAND2_X1 U296 ( .A1(\mem[0][3] ), .A2(n20), .ZN(n24) );
  OAI21_X1 U297 ( .B1(n374), .B2(n393), .A(n36), .ZN(n173) );
  NAND2_X1 U298 ( .A1(\mem[0][15] ), .A2(n20), .ZN(n36) );
  MUX2_X1 U299 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n365), .Z(n1) );
  MUX2_X1 U300 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n364), .Z(n2) );
  MUX2_X1 U301 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U302 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n366), .Z(n4) );
  MUX2_X1 U303 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U304 ( .A(n5), .B(n4), .S(n363), .Z(n6) );
  MUX2_X1 U305 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U306 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U307 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U308 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U309 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U310 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U311 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U312 ( .A(n12), .B(n9), .S(N12), .Z(N27) );
  MUX2_X1 U313 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U314 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U315 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U316 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U317 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U318 ( .A(n17), .B(n16), .S(n363), .Z(n18) );
  MUX2_X1 U319 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U320 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U321 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U322 ( .A(n286), .B(n19), .S(N11), .Z(n287) );
  MUX2_X1 U323 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U324 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U325 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U326 ( .A(n290), .B(n287), .S(N12), .Z(N25) );
  MUX2_X1 U327 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U328 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n366), .Z(n292) );
  MUX2_X1 U329 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U330 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n365), .Z(n294) );
  MUX2_X1 U331 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n364), .Z(n295) );
  MUX2_X1 U332 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U333 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U334 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n366), .Z(n297) );
  MUX2_X1 U335 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n364), .Z(n298) );
  MUX2_X1 U336 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U337 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n366), .Z(n300) );
  MUX2_X1 U338 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U339 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U340 ( .A(n302), .B(n299), .S(N12), .Z(N23) );
  MUX2_X1 U341 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n364), .Z(n303) );
  MUX2_X1 U342 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U343 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U344 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n364), .Z(n306) );
  MUX2_X1 U345 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n366), .Z(n307) );
  MUX2_X1 U346 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U347 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U348 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n365), .Z(n309) );
  MUX2_X1 U349 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n364), .Z(n310) );
  MUX2_X1 U350 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U351 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n365), .Z(n312) );
  MUX2_X1 U352 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n366), .Z(n313) );
  MUX2_X1 U353 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U354 ( .A(n314), .B(n311), .S(N12), .Z(N21) );
  MUX2_X1 U355 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n366), .Z(n315) );
  MUX2_X1 U356 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n316) );
  MUX2_X1 U357 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U358 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n365), .Z(n318) );
  MUX2_X1 U359 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n364), .Z(n319) );
  MUX2_X1 U360 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U361 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U362 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n364), .Z(n321) );
  MUX2_X1 U363 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n365), .Z(n322) );
  MUX2_X1 U364 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U365 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U366 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n364), .Z(n325) );
  MUX2_X1 U367 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U368 ( .A(n326), .B(n323), .S(N12), .Z(N19) );
  MUX2_X1 U369 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n365), .Z(n327) );
  MUX2_X1 U370 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U371 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U372 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n365), .Z(n330) );
  MUX2_X1 U373 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U374 ( .A(n331), .B(n330), .S(N11), .Z(n332) );
  MUX2_X1 U375 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U376 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U377 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U378 ( .A(n334), .B(n333), .S(n363), .Z(n335) );
  MUX2_X1 U379 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U380 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U381 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U382 ( .A(n338), .B(n335), .S(N12), .Z(N17) );
  MUX2_X1 U383 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U384 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U385 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U386 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U387 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U388 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U389 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U390 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U391 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U392 ( .A(n346), .B(n345), .S(n363), .Z(n347) );
  MUX2_X1 U393 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U394 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U395 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U396 ( .A(n350), .B(n347), .S(N12), .Z(N15) );
  MUX2_X1 U397 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U398 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U399 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U400 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U401 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U402 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U403 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U404 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U405 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U406 ( .A(n358), .B(n357), .S(n363), .Z(n359) );
  MUX2_X1 U407 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U408 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U409 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U410 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
  INV_X1 U411 ( .A(data_in[0]), .ZN(n378) );
endmodule


module datapath_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n19, n21, n22, n23, n24, n25, n27, n29, n30, n31, n32, n33, n35, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n51, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70,
         n71, n73, n75, n77, n79, n81, n82, n83, n84, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n155,
         n156;

  FA_X1 U3 ( .A(A[14]), .B(B[14]), .CI(n71), .CO(n16), .S(SUM[14]) );
  OR2_X1 U104 ( .A1(A[0]), .A2(B[0]), .ZN(n140) );
  CLKBUF_X1 U105 ( .A(n22), .Z(n141) );
  CLKBUF_X1 U106 ( .A(n30), .Z(n142) );
  CLKBUF_X1 U107 ( .A(n57), .Z(n143) );
  CLKBUF_X1 U108 ( .A(n41), .Z(n144) );
  CLKBUF_X1 U109 ( .A(n33), .Z(n145) );
  CLKBUF_X1 U110 ( .A(n54), .Z(n146) );
  AOI21_X1 U111 ( .B1(n54), .B2(n153), .A(n51), .ZN(n147) );
  AOI21_X1 U112 ( .B1(n30), .B2(n155), .A(n27), .ZN(n148) );
  NOR2_X1 U113 ( .A1(A[3]), .A2(B[3]), .ZN(n149) );
  INV_X1 U114 ( .A(n37), .ZN(n35) );
  INV_X1 U115 ( .A(n29), .ZN(n27) );
  INV_X1 U116 ( .A(n53), .ZN(n51) );
  INV_X1 U117 ( .A(n45), .ZN(n43) );
  NAND2_X1 U118 ( .A1(n84), .A2(n68), .ZN(n14) );
  INV_X1 U119 ( .A(n67), .ZN(n84) );
  NAND2_X1 U120 ( .A1(n75), .A2(n32), .ZN(n5) );
  INV_X1 U121 ( .A(n31), .ZN(n75) );
  XOR2_X1 U122 ( .A(n65), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U123 ( .A1(n83), .A2(n64), .ZN(n13) );
  AND2_X1 U124 ( .A1(n140), .A2(n70), .ZN(SUM[0]) );
  NAND2_X1 U125 ( .A1(n81), .A2(n56), .ZN(n11) );
  INV_X1 U126 ( .A(n55), .ZN(n81) );
  NAND2_X1 U127 ( .A1(n73), .A2(n24), .ZN(n3) );
  INV_X1 U128 ( .A(n23), .ZN(n73) );
  NAND2_X1 U129 ( .A1(n77), .A2(n40), .ZN(n7) );
  INV_X1 U130 ( .A(n39), .ZN(n77) );
  NAND2_X1 U131 ( .A1(n79), .A2(n48), .ZN(n9) );
  INV_X1 U132 ( .A(n47), .ZN(n79) );
  NAND2_X1 U133 ( .A1(n154), .A2(n21), .ZN(n2) );
  NAND2_X1 U134 ( .A1(n152), .A2(n37), .ZN(n6) );
  NAND2_X1 U135 ( .A1(n151), .A2(n45), .ZN(n8) );
  NAND2_X1 U136 ( .A1(n153), .A2(n53), .ZN(n10) );
  XNOR2_X1 U137 ( .A(n62), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U138 ( .A1(n82), .A2(n61), .ZN(n12) );
  XNOR2_X1 U139 ( .A(n142), .B(n4), .ZN(SUM[11]) );
  NAND2_X1 U140 ( .A1(n155), .A2(n29), .ZN(n4) );
  NOR2_X1 U141 ( .A1(A[3]), .A2(B[3]), .ZN(n60) );
  NOR2_X1 U142 ( .A1(A[1]), .A2(B[1]), .ZN(n67) );
  NAND2_X1 U143 ( .A1(A[2]), .A2(B[2]), .ZN(n64) );
  INV_X1 U144 ( .A(n21), .ZN(n19) );
  NOR2_X1 U145 ( .A1(A[8]), .A2(B[8]), .ZN(n39) );
  NOR2_X1 U146 ( .A1(A[6]), .A2(B[6]), .ZN(n47) );
  NOR2_X1 U147 ( .A1(A[4]), .A2(B[4]), .ZN(n55) );
  NOR2_X1 U148 ( .A1(A[12]), .A2(B[12]), .ZN(n23) );
  NAND2_X1 U149 ( .A1(A[7]), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U150 ( .A1(A[9]), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U151 ( .A1(A[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U152 ( .A1(A[13]), .A2(B[13]), .ZN(n21) );
  NAND2_X1 U153 ( .A1(A[11]), .A2(B[11]), .ZN(n29) );
  NAND2_X1 U154 ( .A1(A[8]), .A2(B[8]), .ZN(n40) );
  NAND2_X1 U155 ( .A1(A[6]), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U156 ( .A1(A[4]), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U157 ( .A1(A[12]), .A2(B[12]), .ZN(n24) );
  OR2_X1 U158 ( .A1(A[7]), .A2(B[7]), .ZN(n151) );
  OR2_X1 U159 ( .A1(A[9]), .A2(B[9]), .ZN(n152) );
  OR2_X1 U160 ( .A1(A[5]), .A2(B[5]), .ZN(n153) );
  OR2_X1 U161 ( .A1(A[13]), .A2(B[13]), .ZN(n154) );
  OR2_X1 U162 ( .A1(A[11]), .A2(B[11]), .ZN(n155) );
  XNOR2_X1 U163 ( .A(n16), .B(n156), .ZN(SUM[15]) );
  XNOR2_X1 U164 ( .A(B[15]), .B(A[15]), .ZN(n156) );
  NAND2_X1 U165 ( .A1(A[10]), .A2(B[10]), .ZN(n32) );
  NOR2_X1 U166 ( .A1(A[10]), .A2(B[10]), .ZN(n31) );
  INV_X1 U167 ( .A(n17), .ZN(n71) );
  OAI21_X1 U168 ( .B1(n33), .B2(n31), .A(n32), .ZN(n30) );
  AOI21_X1 U169 ( .B1(n38), .B2(n152), .A(n35), .ZN(n33) );
  XOR2_X1 U170 ( .A(n14), .B(n70), .Z(SUM[1]) );
  INV_X1 U171 ( .A(n66), .ZN(n65) );
  AOI21_X1 U172 ( .B1(n146), .B2(n153), .A(n51), .ZN(n49) );
  NAND2_X1 U173 ( .A1(A[0]), .A2(B[0]), .ZN(n70) );
  OAI21_X1 U174 ( .B1(n67), .B2(n70), .A(n68), .ZN(n66) );
  OAI21_X1 U175 ( .B1(n57), .B2(n55), .A(n56), .ZN(n54) );
  XNOR2_X1 U176 ( .A(n46), .B(n8), .ZN(SUM[7]) );
  OAI21_X1 U177 ( .B1(n65), .B2(n63), .A(n64), .ZN(n62) );
  INV_X1 U178 ( .A(n63), .ZN(n83) );
  AOI21_X1 U179 ( .B1(n46), .B2(n151), .A(n43), .ZN(n41) );
  NOR2_X1 U180 ( .A1(A[2]), .A2(B[2]), .ZN(n63) );
  OAI21_X1 U181 ( .B1(n147), .B2(n47), .A(n48), .ZN(n46) );
  XOR2_X1 U182 ( .A(n49), .B(n9), .Z(SUM[6]) );
  NAND2_X1 U183 ( .A1(A[1]), .A2(B[1]), .ZN(n68) );
  XNOR2_X1 U184 ( .A(n38), .B(n6), .ZN(SUM[9]) );
  XNOR2_X1 U185 ( .A(n146), .B(n10), .ZN(SUM[5]) );
  XNOR2_X1 U186 ( .A(n141), .B(n2), .ZN(SUM[13]) );
  XOR2_X1 U187 ( .A(n144), .B(n7), .Z(SUM[8]) );
  XOR2_X1 U188 ( .A(n143), .B(n11), .Z(SUM[4]) );
  AOI21_X1 U189 ( .B1(n22), .B2(n154), .A(n19), .ZN(n17) );
  OAI21_X1 U190 ( .B1(n148), .B2(n23), .A(n24), .ZN(n22) );
  OAI21_X1 U191 ( .B1(n41), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U192 ( .B1(n58), .B2(n66), .A(n59), .ZN(n57) );
  AOI21_X1 U193 ( .B1(n142), .B2(n155), .A(n27), .ZN(n25) );
  XOR2_X1 U194 ( .A(n25), .B(n3), .Z(SUM[12]) );
  XOR2_X1 U195 ( .A(n145), .B(n5), .Z(SUM[10]) );
  INV_X1 U196 ( .A(n149), .ZN(n82) );
  NOR2_X1 U197 ( .A1(n63), .A2(n149), .ZN(n58) );
  OAI21_X1 U198 ( .B1(n60), .B2(n64), .A(n61), .ZN(n59) );
  NAND2_X1 U199 ( .A1(A[3]), .A2(B[3]), .ZN(n61) );
endmodule


module datapath_DW_mult_tc_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47,
         n51, n56, n57, n58, n61, n62, n63, n64, n65, n66, n67, n68, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n95, n97, n98, n100, n101, n102, n103, n105,
         n107, n108, n109, n112, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n163, n166, n167, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n248, n249, n250, n251, n253, n254, n255,
         n256, n257, n258, n259, n261, n262, n263, n264, n265, n266, n267,
         n268, n276, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381;
  assign n167 = a[0];
  assign n248 = b[0];
  assign n265 = a[7];
  assign n266 = a[5];
  assign n267 = a[3];
  assign n268 = a[1];

  FA_X1 U131 ( .A(n174), .B(n121), .CI(n181), .CO(n117), .S(n118) );
  FA_X1 U132 ( .A(n122), .B(n175), .CI(n125), .CO(n119), .S(n120) );
  FA_X1 U134 ( .A(n129), .B(n176), .CI(n126), .CO(n123), .S(n124) );
  FA_X1 U135 ( .A(n182), .B(n131), .CI(n189), .CO(n125), .S(n126) );
  FA_X1 U136 ( .A(n135), .B(n137), .CI(n130), .CO(n127), .S(n128) );
  FA_X1 U137 ( .A(n177), .B(n183), .CI(n132), .CO(n129), .S(n130) );
  FA_X1 U140 ( .A(n197), .B(n184), .CI(n143), .CO(n135), .S(n136) );
  FA_X1 U143 ( .A(n147), .B(n144), .CI(n142), .CO(n139), .S(n140) );
  FA_X1 U144 ( .A(n185), .B(n198), .CI(n191), .CO(n141), .S(n142) );
  HA_X1 U145 ( .A(n179), .B(n169), .CO(n143), .S(n144) );
  FA_X1 U146 ( .A(n151), .B(n186), .CI(n148), .CO(n145), .S(n146) );
  FA_X1 U147 ( .A(n199), .B(n180), .CI(n192), .CO(n147), .S(n148) );
  FA_X1 U148 ( .A(n193), .B(n200), .CI(n152), .CO(n149), .S(n150) );
  HA_X1 U149 ( .A(n170), .B(n187), .CO(n151), .S(n152) );
  FA_X1 U150 ( .A(n201), .B(n188), .CI(n194), .CO(n153), .S(n154) );
  HA_X1 U151 ( .A(n195), .B(n202), .CO(n155), .S(n156) );
  OR2_X1 U271 ( .A1(n370), .A2(n167), .ZN(n340) );
  BUF_X2 U272 ( .A(n257), .Z(n379) );
  NOR2_X1 U273 ( .A1(n124), .A2(n127), .ZN(n332) );
  NOR2_X1 U274 ( .A1(n119), .A2(n118), .ZN(n41) );
  INV_X1 U275 ( .A(n317), .ZN(n85) );
  OR2_X1 U276 ( .A1(n120), .A2(n123), .ZN(n306) );
  OR2_X1 U277 ( .A1(n203), .A2(n196), .ZN(n307) );
  OR2_X1 U278 ( .A1(n204), .A2(n172), .ZN(n308) );
  NAND2_X1 U279 ( .A1(n314), .A2(n315), .ZN(n309) );
  CLKBUF_X1 U280 ( .A(n372), .Z(n310) );
  XOR2_X1 U281 ( .A(n264), .B(b[6]), .Z(n233) );
  INV_X1 U282 ( .A(n312), .ZN(n311) );
  CLKBUF_X1 U283 ( .A(n266), .Z(n344) );
  NAND2_X1 U284 ( .A1(n266), .A2(n313), .ZN(n314) );
  NAND2_X1 U285 ( .A1(n312), .A2(a[4]), .ZN(n315) );
  NAND2_X1 U286 ( .A1(n314), .A2(n315), .ZN(n250) );
  INV_X1 U287 ( .A(n266), .ZN(n312) );
  INV_X1 U288 ( .A(a[4]), .ZN(n313) );
  BUF_X1 U289 ( .A(n267), .Z(n381) );
  CLKBUF_X1 U290 ( .A(n268), .Z(n316) );
  OR2_X1 U291 ( .A1(n370), .A2(n167), .ZN(n256) );
  OR2_X1 U292 ( .A1(n370), .A2(n167), .ZN(n341) );
  OAI22_X1 U293 ( .A1(n375), .A2(n224), .B1(n223), .B2(n259), .ZN(n131) );
  AND2_X2 U294 ( .A1(n150), .A2(n153), .ZN(n317) );
  CLKBUF_X1 U295 ( .A(n80), .Z(n318) );
  NOR2_X1 U296 ( .A1(n146), .A2(n149), .ZN(n319) );
  AND2_X1 U297 ( .A1(n306), .A2(n103), .ZN(n39) );
  NOR2_X1 U298 ( .A1(n41), .A2(n34), .ZN(n320) );
  CLKBUF_X1 U299 ( .A(n255), .Z(n321) );
  XNOR2_X1 U300 ( .A(n136), .B(n338), .ZN(n322) );
  NAND2_X1 U301 ( .A1(n357), .A2(a[2]), .ZN(n323) );
  OR2_X1 U302 ( .A1(n154), .A2(n155), .ZN(n324) );
  CLKBUF_X1 U303 ( .A(n330), .Z(n325) );
  NOR2_X1 U304 ( .A1(n66), .A2(n61), .ZN(n326) );
  NOR2_X1 U305 ( .A1(n66), .A2(n61), .ZN(n3) );
  AND2_X1 U306 ( .A1(n120), .A2(n123), .ZN(n327) );
  NOR2_X1 U307 ( .A1(n146), .A2(n149), .ZN(n79) );
  CLKBUF_X1 U308 ( .A(n306), .Z(n328) );
  CLKBUF_X1 U309 ( .A(n331), .Z(n329) );
  OAI21_X1 U310 ( .B1(n332), .B2(n67), .A(n62), .ZN(n330) );
  OAI21_X1 U311 ( .B1(n67), .B2(n332), .A(n62), .ZN(n2) );
  OAI21_X2 U312 ( .B1(n87), .B2(n89), .A(n88), .ZN(n86) );
  AOI21_X1 U313 ( .B1(n363), .B2(n353), .A(n336), .ZN(n331) );
  AOI21_X1 U314 ( .B1(n363), .B2(n353), .A(n336), .ZN(n366) );
  NOR2_X1 U315 ( .A1(n124), .A2(n127), .ZN(n61) );
  NAND2_X2 U316 ( .A1(n249), .A2(n337), .ZN(n253) );
  CLKBUF_X1 U317 ( .A(n268), .Z(n333) );
  XOR2_X1 U318 ( .A(n268), .B(a[2]), .Z(n334) );
  NAND2_X1 U319 ( .A1(n360), .A2(n359), .ZN(n335) );
  OAI21_X1 U320 ( .B1(n76), .B2(n72), .A(n73), .ZN(n336) );
  XNOR2_X1 U321 ( .A(n266), .B(a[6]), .ZN(n337) );
  XNOR2_X1 U322 ( .A(n136), .B(n338), .ZN(n134) );
  XNOR2_X1 U323 ( .A(n141), .B(n138), .ZN(n338) );
  XNOR2_X1 U324 ( .A(n190), .B(n178), .ZN(n138) );
  CLKBUF_X1 U325 ( .A(n377), .Z(n339) );
  CLKBUF_X1 U326 ( .A(n75), .Z(n342) );
  XNOR2_X1 U327 ( .A(n351), .B(a[4]), .ZN(n343) );
  CLKBUF_X3 U328 ( .A(n267), .Z(n351) );
  CLKBUF_X1 U329 ( .A(n266), .Z(n369) );
  NAND2_X1 U330 ( .A1(n136), .A2(n141), .ZN(n345) );
  NAND2_X1 U331 ( .A1(n136), .A2(n138), .ZN(n346) );
  NAND2_X1 U332 ( .A1(n141), .A2(n138), .ZN(n347) );
  NAND3_X1 U333 ( .A1(n345), .A2(n346), .A3(n347), .ZN(n133) );
  AOI21_X1 U334 ( .B1(n368), .B2(n86), .A(n317), .ZN(n348) );
  XNOR2_X1 U335 ( .A(n63), .B(n349), .ZN(product[10]) );
  AND2_X1 U336 ( .A1(n105), .A2(n62), .ZN(n349) );
  CLKBUF_X1 U337 ( .A(n267), .Z(n350) );
  CLKBUF_X1 U338 ( .A(n76), .Z(n352) );
  NOR2_X1 U339 ( .A1(n377), .A2(n75), .ZN(n353) );
  INV_X1 U340 ( .A(n334), .ZN(n354) );
  XNOR2_X1 U341 ( .A(n268), .B(a[2]), .ZN(n259) );
  XNOR2_X1 U342 ( .A(n268), .B(a[2]), .ZN(n362) );
  AOI21_X1 U343 ( .B1(n368), .B2(n86), .A(n317), .ZN(n355) );
  AOI21_X1 U344 ( .B1(n368), .B2(n86), .A(n317), .ZN(n81) );
  AOI21_X1 U345 ( .B1(n320), .B2(n327), .A(n33), .ZN(n356) );
  NAND2_X1 U346 ( .A1(n351), .A2(n358), .ZN(n359) );
  NAND2_X1 U347 ( .A1(n357), .A2(a[2]), .ZN(n360) );
  NAND2_X1 U348 ( .A1(n323), .A2(n359), .ZN(n251) );
  INV_X1 U349 ( .A(n381), .ZN(n357) );
  INV_X1 U350 ( .A(a[2]), .ZN(n358) );
  INV_X1 U351 ( .A(n65), .ZN(n361) );
  BUF_X2 U352 ( .A(n265), .Z(n378) );
  OAI21_X1 U353 ( .B1(n355), .B2(n79), .A(n80), .ZN(n363) );
  OAI21_X1 U354 ( .B1(n319), .B2(n348), .A(n80), .ZN(n364) );
  CLKBUF_X1 U355 ( .A(n3), .Z(n365) );
  NOR2_X1 U356 ( .A1(n117), .A2(n116), .ZN(n34) );
  AOI21_X1 U357 ( .B1(n78), .B2(n70), .A(n71), .ZN(n1) );
  INV_X1 U358 ( .A(n66), .ZN(n64) );
  INV_X1 U359 ( .A(n67), .ZN(n65) );
  OAI21_X1 U360 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NOR2_X1 U361 ( .A1(n41), .A2(n34), .ZN(n32) );
  INV_X1 U362 ( .A(n23), .ZN(n101) );
  INV_X1 U363 ( .A(n34), .ZN(n102) );
  NOR2_X1 U364 ( .A1(n140), .A2(n145), .ZN(n75) );
  INV_X1 U365 ( .A(n115), .ZN(n116) );
  NAND2_X1 U366 ( .A1(n119), .A2(n118), .ZN(n44) );
  NAND2_X1 U367 ( .A1(n140), .A2(n145), .ZN(n76) );
  AOI21_X1 U368 ( .B1(n307), .B2(n98), .A(n95), .ZN(n93) );
  INV_X1 U369 ( .A(n97), .ZN(n95) );
  NOR2_X1 U370 ( .A1(n173), .A2(n115), .ZN(n23) );
  NAND2_X1 U371 ( .A1(n173), .A2(n115), .ZN(n24) );
  INV_X1 U372 ( .A(n100), .ZN(n98) );
  NAND2_X1 U373 ( .A1(n117), .A2(n116), .ZN(n35) );
  NAND2_X1 U374 ( .A1(n124), .A2(n127), .ZN(n62) );
  NAND2_X1 U375 ( .A1(n120), .A2(n123), .ZN(n51) );
  NAND2_X1 U376 ( .A1(n64), .A2(n361), .ZN(n9) );
  NAND2_X1 U377 ( .A1(n109), .A2(n318), .ZN(n12) );
  INV_X1 U378 ( .A(n319), .ZN(n109) );
  XOR2_X1 U379 ( .A(n15), .B(n93), .Z(product[3]) );
  INV_X1 U380 ( .A(n91), .ZN(n112) );
  XOR2_X1 U381 ( .A(n14), .B(n89), .Z(product[4]) );
  NAND2_X1 U382 ( .A1(n324), .A2(n88), .ZN(n14) );
  XOR2_X1 U383 ( .A(n77), .B(n11), .Z(product[7]) );
  NAND2_X1 U384 ( .A1(n108), .A2(n352), .ZN(n11) );
  INV_X1 U385 ( .A(n342), .ZN(n108) );
  NAND2_X1 U386 ( .A1(n101), .A2(n24), .ZN(n4) );
  OAI21_X1 U387 ( .B1(n77), .B2(n342), .A(n352), .ZN(n74) );
  XNOR2_X1 U388 ( .A(n45), .B(n6), .ZN(product[12]) );
  NAND2_X1 U389 ( .A1(n103), .A2(n44), .ZN(n6) );
  XNOR2_X1 U390 ( .A(n36), .B(n5), .ZN(product[13]) );
  NAND2_X1 U391 ( .A1(n102), .A2(n35), .ZN(n5) );
  XNOR2_X1 U392 ( .A(n56), .B(n7), .ZN(product[11]) );
  XNOR2_X1 U393 ( .A(n16), .B(n98), .ZN(product[2]) );
  NAND2_X1 U394 ( .A1(n307), .A2(n97), .ZN(n16) );
  AND2_X1 U395 ( .A1(n308), .A2(n100), .ZN(product[1]) );
  INV_X1 U396 ( .A(n160), .ZN(n181) );
  INV_X1 U397 ( .A(n121), .ZN(n122) );
  NOR2_X1 U398 ( .A1(n154), .A2(n155), .ZN(n87) );
  INV_X1 U399 ( .A(n157), .ZN(n173) );
  OR2_X1 U400 ( .A1(n150), .A2(n153), .ZN(n368) );
  OR2_X1 U401 ( .A1(n248), .A2(n263), .ZN(n231) );
  XNOR2_X1 U402 ( .A(n378), .B(b[7]), .ZN(n205) );
  XNOR2_X1 U403 ( .A(n378), .B(b[4]), .ZN(n208) );
  XNOR2_X1 U404 ( .A(n378), .B(b[6]), .ZN(n206) );
  XNOR2_X1 U405 ( .A(n378), .B(b[3]), .ZN(n209) );
  XNOR2_X1 U406 ( .A(n378), .B(b[5]), .ZN(n207) );
  XNOR2_X1 U407 ( .A(n378), .B(b[1]), .ZN(n211) );
  XNOR2_X1 U408 ( .A(n378), .B(b[2]), .ZN(n210) );
  XNOR2_X1 U409 ( .A(n378), .B(n248), .ZN(n212) );
  AND2_X1 U410 ( .A1(n248), .A2(n161), .ZN(n188) );
  AND2_X1 U411 ( .A1(n248), .A2(n158), .ZN(n180) );
  OR2_X1 U412 ( .A1(n248), .A2(n261), .ZN(n213) );
  INV_X1 U413 ( .A(n265), .ZN(n261) );
  OR2_X1 U414 ( .A1(n248), .A2(n262), .ZN(n222) );
  AND2_X1 U415 ( .A1(n248), .A2(n167), .ZN(product[0]) );
  INV_X1 U416 ( .A(n332), .ZN(n105) );
  NOR2_X1 U417 ( .A1(n30), .A2(n23), .ZN(n21) );
  INV_X1 U418 ( .A(n30), .ZN(n28) );
  NAND2_X1 U419 ( .A1(n368), .A2(n85), .ZN(n13) );
  XNOR2_X1 U420 ( .A(n13), .B(n86), .ZN(product[5]) );
  XNOR2_X1 U421 ( .A(n268), .B(n167), .ZN(n370) );
  INV_X1 U422 ( .A(n167), .ZN(n276) );
  NAND2_X1 U423 ( .A1(n258), .A2(n309), .ZN(n371) );
  NAND2_X1 U424 ( .A1(n250), .A2(n380), .ZN(n372) );
  NAND2_X1 U425 ( .A1(n258), .A2(n309), .ZN(n254) );
  BUF_X1 U426 ( .A(n258), .Z(n373) );
  NAND2_X1 U427 ( .A1(n335), .A2(n259), .ZN(n374) );
  NAND2_X1 U428 ( .A1(n362), .A2(n251), .ZN(n375) );
  NAND2_X1 U429 ( .A1(n335), .A2(n362), .ZN(n255) );
  OR2_X1 U430 ( .A1(n248), .A2(n264), .ZN(n240) );
  OR2_X1 U431 ( .A1(n190), .A2(n178), .ZN(n137) );
  AND2_X1 U432 ( .A1(n248), .A2(n334), .ZN(n196) );
  INV_X1 U433 ( .A(n166), .ZN(n197) );
  CLKBUF_X1 U434 ( .A(n68), .Z(n376) );
  XNOR2_X1 U435 ( .A(n376), .B(n9), .ZN(product[9]) );
  XNOR2_X1 U436 ( .A(n74), .B(n10), .ZN(product[8]) );
  INV_X1 U437 ( .A(n90), .ZN(n89) );
  NAND2_X1 U438 ( .A1(n154), .A2(n155), .ZN(n88) );
  NAND2_X1 U439 ( .A1(n107), .A2(n73), .ZN(n10) );
  NAND2_X1 U440 ( .A1(n322), .A2(n139), .ZN(n73) );
  NAND2_X1 U441 ( .A1(n146), .A2(n149), .ZN(n80) );
  INV_X1 U442 ( .A(n330), .ZN(n58) );
  NOR2_X1 U443 ( .A1(n133), .A2(n128), .ZN(n66) );
  NAND2_X1 U444 ( .A1(n128), .A2(n133), .ZN(n67) );
  NOR2_X1 U445 ( .A1(n322), .A2(n139), .ZN(n377) );
  NOR2_X1 U446 ( .A1(n134), .A2(n139), .ZN(n72) );
  XNOR2_X1 U447 ( .A(n266), .B(a[6]), .ZN(n257) );
  OAI21_X1 U448 ( .B1(n91), .B2(n93), .A(n92), .ZN(n90) );
  NAND2_X1 U449 ( .A1(n112), .A2(n92), .ZN(n15) );
  INV_X1 U450 ( .A(n163), .ZN(n189) );
  XNOR2_X1 U451 ( .A(n351), .B(a[4]), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(a[4]), .ZN(n258) );
  XOR2_X1 U453 ( .A(n265), .B(a[6]), .Z(n249) );
  INV_X1 U454 ( .A(n31), .ZN(n29) );
  OAI21_X1 U455 ( .B1(n356), .B2(n23), .A(n24), .ZN(n22) );
  AOI21_X1 U456 ( .B1(n32), .B2(n327), .A(n33), .ZN(n31) );
  XNOR2_X1 U457 ( .A(n25), .B(n4), .ZN(product[14]) );
  NAND2_X1 U458 ( .A1(n203), .A2(n196), .ZN(n97) );
  INV_X1 U459 ( .A(n18), .ZN(product[15]) );
  AOI21_X1 U460 ( .B1(n325), .B2(n21), .A(n22), .ZN(n20) );
  OAI22_X1 U461 ( .A1(n341), .A2(n235), .B1(n234), .B2(n276), .ZN(n200) );
  OAI22_X1 U462 ( .A1(n340), .A2(n236), .B1(n235), .B2(n276), .ZN(n201) );
  NAND2_X1 U463 ( .A1(n204), .A2(n172), .ZN(n100) );
  OAI22_X1 U464 ( .A1(n341), .A2(n234), .B1(n233), .B2(n276), .ZN(n199) );
  OAI22_X1 U465 ( .A1(n256), .A2(n233), .B1(n232), .B2(n276), .ZN(n198) );
  OAI22_X1 U466 ( .A1(n232), .A2(n340), .B1(n232), .B2(n276), .ZN(n166) );
  OAI22_X1 U467 ( .A1(n340), .A2(n237), .B1(n236), .B2(n276), .ZN(n202) );
  OAI22_X1 U468 ( .A1(n256), .A2(n238), .B1(n237), .B2(n276), .ZN(n203) );
  OAI22_X1 U469 ( .A1(n256), .A2(n239), .B1(n238), .B2(n276), .ZN(n204) );
  OAI22_X1 U470 ( .A1(n341), .A2(n264), .B1(n240), .B2(n276), .ZN(n172) );
  INV_X1 U471 ( .A(n131), .ZN(n132) );
  AOI21_X1 U472 ( .B1(n2), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U473 ( .B1(n330), .B2(n28), .A(n29), .ZN(n27) );
  NAND2_X1 U474 ( .A1(n156), .A2(n171), .ZN(n92) );
  NOR2_X1 U475 ( .A1(n156), .A2(n171), .ZN(n91) );
  NAND2_X1 U476 ( .A1(n3), .A2(n28), .ZN(n26) );
  NAND2_X1 U477 ( .A1(n39), .A2(n3), .ZN(n37) );
  INV_X1 U478 ( .A(n326), .ZN(n57) );
  NAND2_X1 U479 ( .A1(n365), .A2(n21), .ZN(n19) );
  INV_X1 U480 ( .A(n339), .ZN(n107) );
  NOR2_X1 U481 ( .A1(n75), .A2(n377), .ZN(n70) );
  OAI21_X1 U482 ( .B1(n72), .B2(n76), .A(n73), .ZN(n71) );
  OAI22_X1 U483 ( .A1(n371), .A2(n220), .B1(n343), .B2(n219), .ZN(n186) );
  OAI22_X1 U484 ( .A1(n310), .A2(n215), .B1(n373), .B2(n214), .ZN(n121) );
  INV_X1 U485 ( .A(n373), .ZN(n161) );
  OAI22_X1 U486 ( .A1(n214), .A2(n310), .B1(n214), .B2(n343), .ZN(n160) );
  OAI22_X1 U487 ( .A1(n372), .A2(n219), .B1(n373), .B2(n218), .ZN(n185) );
  OAI22_X1 U488 ( .A1(n372), .A2(n218), .B1(n373), .B2(n217), .ZN(n184) );
  OAI22_X1 U489 ( .A1(n371), .A2(n217), .B1(n343), .B2(n216), .ZN(n183) );
  OAI22_X1 U490 ( .A1(n371), .A2(n216), .B1(n343), .B2(n215), .ZN(n182) );
  XNOR2_X1 U491 ( .A(n351), .B(b[2]), .ZN(n228) );
  OAI22_X1 U492 ( .A1(n254), .A2(n262), .B1(n222), .B2(n343), .ZN(n170) );
  OAI22_X1 U493 ( .A1(n254), .A2(n221), .B1(n220), .B2(n380), .ZN(n187) );
  XNOR2_X1 U494 ( .A(n350), .B(b[3]), .ZN(n227) );
  XNOR2_X1 U495 ( .A(n351), .B(b[4]), .ZN(n226) );
  INV_X1 U496 ( .A(n350), .ZN(n263) );
  XNOR2_X1 U497 ( .A(n350), .B(b[5]), .ZN(n225) );
  XNOR2_X1 U498 ( .A(n351), .B(b[6]), .ZN(n224) );
  XNOR2_X1 U499 ( .A(n350), .B(n248), .ZN(n230) );
  XNOR2_X1 U500 ( .A(n350), .B(b[7]), .ZN(n223) );
  XNOR2_X1 U501 ( .A(n351), .B(b[1]), .ZN(n229) );
  INV_X1 U502 ( .A(n41), .ZN(n103) );
  OAI21_X1 U503 ( .B1(n51), .B2(n41), .A(n44), .ZN(n40) );
  OAI22_X1 U504 ( .A1(n374), .A2(n228), .B1(n259), .B2(n227), .ZN(n193) );
  OAI22_X1 U505 ( .A1(n374), .A2(n229), .B1(n354), .B2(n228), .ZN(n194) );
  OAI22_X1 U506 ( .A1(n321), .A2(n263), .B1(n231), .B2(n354), .ZN(n171) );
  OAI22_X1 U507 ( .A1(n374), .A2(n225), .B1(n354), .B2(n224), .ZN(n190) );
  OAI22_X1 U508 ( .A1(n255), .A2(n227), .B1(n259), .B2(n226), .ZN(n192) );
  OAI22_X1 U509 ( .A1(n255), .A2(n226), .B1(n259), .B2(n225), .ZN(n191) );
  XNOR2_X1 U510 ( .A(n316), .B(b[4]), .ZN(n235) );
  XNOR2_X1 U511 ( .A(n316), .B(b[5]), .ZN(n234) );
  OAI22_X1 U512 ( .A1(n230), .A2(n255), .B1(n354), .B2(n229), .ZN(n195) );
  OAI22_X1 U513 ( .A1(n223), .A2(n375), .B1(n223), .B2(n259), .ZN(n163) );
  XNOR2_X1 U514 ( .A(n333), .B(b[3]), .ZN(n236) );
  XNOR2_X1 U515 ( .A(n333), .B(b[2]), .ZN(n237) );
  XNOR2_X1 U516 ( .A(n333), .B(n248), .ZN(n239) );
  XNOR2_X1 U517 ( .A(n268), .B(b[7]), .ZN(n232) );
  XNOR2_X1 U518 ( .A(n316), .B(b[1]), .ZN(n238) );
  INV_X1 U519 ( .A(n268), .ZN(n264) );
  INV_X1 U520 ( .A(n364), .ZN(n77) );
  OAI21_X1 U521 ( .B1(n79), .B2(n81), .A(n80), .ZN(n78) );
  XOR2_X1 U522 ( .A(n12), .B(n348), .Z(product[6]) );
  OAI22_X1 U523 ( .A1(n205), .A2(n253), .B1(n205), .B2(n379), .ZN(n157) );
  OAI22_X1 U524 ( .A1(n253), .A2(n209), .B1(n379), .B2(n208), .ZN(n176) );
  OAI22_X1 U525 ( .A1(n253), .A2(n208), .B1(n379), .B2(n207), .ZN(n175) );
  OAI22_X1 U526 ( .A1(n253), .A2(n206), .B1(n379), .B2(n205), .ZN(n115) );
  OAI22_X1 U527 ( .A1(n253), .A2(n207), .B1(n379), .B2(n206), .ZN(n174) );
  INV_X1 U528 ( .A(n379), .ZN(n158) );
  OAI22_X1 U529 ( .A1(n253), .A2(n211), .B1(n379), .B2(n210), .ZN(n178) );
  OAI22_X1 U530 ( .A1(n253), .A2(n210), .B1(n379), .B2(n209), .ZN(n177) );
  OAI22_X1 U531 ( .A1(n253), .A2(n261), .B1(n213), .B2(n379), .ZN(n169) );
  OAI22_X1 U532 ( .A1(n253), .A2(n212), .B1(n379), .B2(n211), .ZN(n179) );
  XNOR2_X1 U533 ( .A(n311), .B(b[2]), .ZN(n219) );
  XNOR2_X1 U534 ( .A(n344), .B(b[5]), .ZN(n216) );
  XNOR2_X1 U535 ( .A(n344), .B(b[6]), .ZN(n215) );
  XNOR2_X1 U536 ( .A(n311), .B(b[7]), .ZN(n214) );
  XNOR2_X1 U537 ( .A(n344), .B(b[3]), .ZN(n218) );
  XNOR2_X1 U538 ( .A(n311), .B(b[4]), .ZN(n217) );
  XNOR2_X1 U539 ( .A(n311), .B(n248), .ZN(n221) );
  INV_X1 U540 ( .A(n369), .ZN(n262) );
  XNOR2_X1 U541 ( .A(n369), .B(b[1]), .ZN(n220) );
  AOI21_X1 U542 ( .B1(n2), .B2(n328), .A(n327), .ZN(n47) );
  NAND2_X1 U543 ( .A1(n326), .A2(n328), .ZN(n46) );
  NAND2_X1 U544 ( .A1(n328), .A2(n51), .ZN(n7) );
  NAND2_X1 U545 ( .A1(n306), .A2(n320), .ZN(n30) );
  OAI21_X1 U546 ( .B1(n329), .B2(n19), .A(n20), .ZN(n18) );
  INV_X1 U547 ( .A(n1), .ZN(n68) );
  OAI21_X1 U548 ( .B1(n366), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U549 ( .B1(n331), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U550 ( .B1(n331), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U551 ( .B1(n366), .B2(n26), .A(n27), .ZN(n25) );
  AOI21_X1 U552 ( .B1(n68), .B2(n64), .A(n65), .ZN(n63) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a, wr_en_a, addr_y, 
        wr_en_y, clear_acc, data_out );
  input [7:0] data_in;
  input [2:0] addr_x;
  input [5:0] addr_a;
  input [2:0] addr_y;
  output [15:0] data_out;
  input clk, wr_en_x, wr_en_a, wr_en_y, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, n2, n3, n4;
  wire   [7:0] data_out_x;
  wire   [7:0] data_out_a;
  wire   [15:0] f;
  wire   [15:0] mul_out_r;
  wire   [15:0] add_r;
  wire   [15:0] mul_out;

  DFF_X1 \mul_out_r_reg[15]  ( .D(N34), .CK(clk), .Q(mul_out_r[15]) );
  DFF_X1 \mul_out_r_reg[14]  ( .D(N33), .CK(clk), .Q(mul_out_r[14]) );
  DFF_X1 \mul_out_r_reg[11]  ( .D(N30), .CK(clk), .Q(mul_out_r[11]) );
  DFF_X1 \mul_out_r_reg[9]  ( .D(N28), .CK(clk), .Q(mul_out_r[9]) );
  DFF_X1 \mul_out_r_reg[8]  ( .D(N27), .CK(clk), .Q(mul_out_r[8]) );
  DFF_X1 \mul_out_r_reg[7]  ( .D(N26), .CK(clk), .Q(mul_out_r[7]) );
  DFF_X1 \mul_out_r_reg[6]  ( .D(N25), .CK(clk), .Q(mul_out_r[6]) );
  DFF_X1 \mul_out_r_reg[5]  ( .D(N24), .CK(clk), .Q(mul_out_r[5]) );
  DFF_X1 \mul_out_r_reg[4]  ( .D(N23), .CK(clk), .Q(mul_out_r[4]) );
  DFF_X1 \mul_out_r_reg[3]  ( .D(N22), .CK(clk), .Q(mul_out_r[3]) );
  DFF_X1 \mul_out_r_reg[2]  ( .D(N21), .CK(clk), .Q(mul_out_r[2]) );
  DFF_X1 \mul_out_r_reg[1]  ( .D(N20), .CK(clk), .Q(mul_out_r[1]) );
  DFF_X1 \mul_out_r_reg[0]  ( .D(N19), .CK(clk), .Q(mul_out_r[0]) );
  DFF_X1 \f_reg[0]  ( .D(N3), .CK(clk), .Q(f[0]) );
  DFF_X1 \f_reg[1]  ( .D(N4), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[2]  ( .D(N5), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(N6), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(N7), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(N8), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[6]  ( .D(N9), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(N10), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[8]  ( .D(N11), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[9]  ( .D(N12), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[10]  ( .D(N13), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[11]  ( .D(N14), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg[12]  ( .D(N15), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[13]  ( .D(N16), .CK(clk), .Q(f[13]) );
  DFF_X1 \f_reg[14]  ( .D(N17), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[15]  ( .D(N18), .CK(clk), .Q(f[15]) );
  memory_WIDTH8_SIZE8_LOGSIZE3 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE64_LOGSIZE6 mem_a ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a), .addr(addr_a), .wr_en(wr_en_a) );
  memory_WIDTH16_SIZE8_LOGSIZE3 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW01_add_1 add_68 ( .A(f), .B(mul_out_r), .CI(1'b0), .SUM(add_r) );
  datapath_DW_mult_tc_1 mult_67 ( .a(data_out_a), .b(data_out_x), .product(
        mul_out) );
  DFF_X1 \mul_out_r_reg[12]  ( .D(N31), .CK(clk), .Q(mul_out_r[12]) );
  DFF_X1 \mul_out_r_reg[13]  ( .D(N32), .CK(clk), .Q(mul_out_r[13]) );
  DFF_X1 \mul_out_r_reg[10]  ( .D(N29), .CK(clk), .Q(mul_out_r[10]) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(clear_acc), .ZN(n4) );
  AND2_X1 U7 ( .A1(add_r[14]), .A2(n3), .ZN(N17) );
  AND2_X1 U8 ( .A1(add_r[13]), .A2(n3), .ZN(N16) );
  AND2_X1 U9 ( .A1(add_r[12]), .A2(n3), .ZN(N15) );
  AND2_X1 U10 ( .A1(add_r[11]), .A2(n3), .ZN(N14) );
  AND2_X1 U11 ( .A1(add_r[10]), .A2(n3), .ZN(N13) );
  AND2_X1 U12 ( .A1(add_r[9]), .A2(n3), .ZN(N12) );
  AND2_X1 U13 ( .A1(add_r[8]), .A2(n3), .ZN(N11) );
  AND2_X1 U14 ( .A1(add_r[7]), .A2(n3), .ZN(N10) );
  AND2_X1 U15 ( .A1(add_r[6]), .A2(n3), .ZN(N9) );
  AND2_X1 U16 ( .A1(add_r[5]), .A2(n3), .ZN(N8) );
  AND2_X1 U17 ( .A1(add_r[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U18 ( .A1(add_r[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U19 ( .A1(add_r[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U20 ( .A1(add_r[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U21 ( .A1(add_r[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U22 ( .A1(mul_out[15]), .A2(n2), .ZN(N34) );
  AND2_X1 U23 ( .A1(mul_out[14]), .A2(n2), .ZN(N33) );
  AND2_X1 U24 ( .A1(mul_out[13]), .A2(n2), .ZN(N32) );
  AND2_X1 U25 ( .A1(mul_out[12]), .A2(n2), .ZN(N31) );
  AND2_X1 U26 ( .A1(mul_out[11]), .A2(n2), .ZN(N30) );
  AND2_X1 U27 ( .A1(mul_out[10]), .A2(n2), .ZN(N29) );
  AND2_X1 U28 ( .A1(mul_out[9]), .A2(n3), .ZN(N28) );
  AND2_X1 U29 ( .A1(mul_out[8]), .A2(n4), .ZN(N27) );
  AND2_X1 U30 ( .A1(mul_out[7]), .A2(n4), .ZN(N26) );
  AND2_X1 U31 ( .A1(mul_out[6]), .A2(n4), .ZN(N25) );
  AND2_X1 U32 ( .A1(mul_out[5]), .A2(n4), .ZN(N24) );
  AND2_X1 U33 ( .A1(mul_out[4]), .A2(n4), .ZN(N23) );
  AND2_X1 U34 ( .A1(mul_out[3]), .A2(n4), .ZN(N22) );
  AND2_X1 U35 ( .A1(mul_out[2]), .A2(n4), .ZN(N21) );
  AND2_X1 U36 ( .A1(mul_out[1]), .A2(n4), .ZN(N20) );
  AND2_X1 U37 ( .A1(mul_out[0]), .A2(n4), .ZN(N19) );
  AND2_X1 U38 ( .A1(add_r[15]), .A2(n4), .ZN(N18) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a, wr_en_a, 
        clear_acc, addr_y, wr_en_y, done, loadMatrix, loadVector );
  output [2:0] addr_x;
  output [5:0] addr_a;
  output [2:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a, clear_acc, wr_en_y, done;
  wire   N17, N18, N19, N20, N21, N26, N27, N28, N29, N30, N44, N45, N46, N54,
         N55, N56, N59, N66, n39, n40, n41, n42, n44, n46, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, \add_103/carry[5] , \add_103/carry[4] ,
         \add_103/carry[3] , \add_103/carry[2] , n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30;
  wire   [3:0] state;

  DFF_X1 \addr_y_reg[0]  ( .D(N54), .CK(clk), .Q(addr_y[0]) );
  DFF_X1 \addr_y_reg[2]  ( .D(N56), .CK(clk), .Q(addr_y[2]), .QN(n44) );
  DFF_X1 \state_reg[0]  ( .D(N17), .CK(clk), .Q(state[0]), .QN(n41) );
  DFF_X1 \state_reg[1]  ( .D(N18), .CK(clk), .Q(state[1]), .QN(n40) );
  DFF_X1 done_reg ( .D(N21), .CK(clk), .Q(done) );
  DFF_X1 \state_reg[2]  ( .D(N19), .CK(clk), .Q(state[2]), .QN(n39) );
  DFF_X1 \state_reg[3]  ( .D(N20), .CK(clk), .Q(state[3]), .QN(n5) );
  DFF_X1 \addr_y_reg[1]  ( .D(N55), .CK(clk), .Q(addr_y[1]), .QN(n46) );
  DFF_X1 \addr_x_reg[0]  ( .D(N44), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N45), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 \addr_x_reg[2]  ( .D(N46), .CK(clk), .Q(addr_x[2]), .QN(n42) );
  DFF_X1 \addr_a_reg[0]  ( .D(n10), .CK(clk), .Q(addr_a[0]), .QN(n2) );
  DFF_X1 \addr_a_reg[5]  ( .D(n15), .CK(clk), .Q(addr_a[5]) );
  DFF_X1 \addr_a_reg[4]  ( .D(n14), .CK(clk), .Q(addr_a[4]) );
  DFF_X1 \addr_a_reg[3]  ( .D(n13), .CK(clk), .Q(addr_a[3]) );
  DFF_X1 \addr_a_reg[2]  ( .D(n12), .CK(clk), .Q(addr_a[2]) );
  DFF_X1 \addr_a_reg[1]  ( .D(n11), .CK(clk), .Q(addr_a[1]) );
  DFF_X1 clear_acc_reg ( .D(N59), .CK(clk), .Q(clear_acc) );
  NAND3_X1 U82 ( .A1(n25), .A2(n46), .A3(addr_y[0]), .ZN(n51) );
  NAND3_X1 U83 ( .A1(n54), .A2(n52), .A3(addr_y[0]), .ZN(n53) );
  NAND3_X1 U84 ( .A1(addr_x[0]), .A2(n57), .A3(addr_x[1]), .ZN(n56) );
  NAND3_X1 U85 ( .A1(n60), .A2(n16), .A3(n74), .ZN(n63) );
  NAND3_X1 U86 ( .A1(n75), .A2(n76), .A3(N66), .ZN(n74) );
  NAND3_X1 U87 ( .A1(n77), .A2(n73), .A3(n75), .ZN(n60) );
  NAND3_X1 U88 ( .A1(n79), .A2(n71), .A3(n70), .ZN(n78) );
  NAND3_X1 U89 ( .A1(n59), .A2(n72), .A3(n80), .ZN(N59) );
  NAND3_X1 U91 ( .A1(n41), .A2(n40), .A3(n55), .ZN(n71) );
  NAND3_X1 U92 ( .A1(n100), .A2(n39), .A3(state[3]), .ZN(n70) );
  NAND3_X1 U93 ( .A1(addr_y[1]), .A2(addr_y[0]), .A3(addr_y[2]), .ZN(n88) );
  NAND3_X1 U94 ( .A1(n99), .A2(n39), .A3(state[3]), .ZN(n80) );
  NAND3_X1 U95 ( .A1(n41), .A2(n40), .A3(n98), .ZN(n54) );
  NAND3_X1 U96 ( .A1(state[1]), .A2(state[0]), .A3(n98), .ZN(n76) );
  NAND3_X1 U97 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n81) );
  HA_X1 \add_103/U1_1_1  ( .A(addr_a[1]), .B(addr_a[0]), .CO(
        \add_103/carry[2] ), .S(N26) );
  HA_X1 \add_103/U1_1_2  ( .A(addr_a[2]), .B(\add_103/carry[2] ), .CO(
        \add_103/carry[3] ), .S(N27) );
  HA_X1 \add_103/U1_1_3  ( .A(addr_a[3]), .B(\add_103/carry[3] ), .CO(
        \add_103/carry[4] ), .S(N28) );
  HA_X1 \add_103/U1_1_4  ( .A(addr_a[4]), .B(\add_103/carry[4] ), .CO(
        \add_103/carry[5] ), .S(N29) );
  INV_X1 U3 ( .A(n57), .ZN(n17) );
  OAI21_X1 U4 ( .B1(n29), .B2(n59), .A(n60), .ZN(n57) );
  NAND2_X1 U5 ( .A1(n29), .A2(n27), .ZN(n73) );
  INV_X1 U6 ( .A(n59), .ZN(n23) );
  INV_X1 U7 ( .A(wr_en_y), .ZN(n16) );
  NOR2_X1 U8 ( .A1(n63), .A2(n69), .ZN(n62) );
  AND4_X1 U9 ( .A1(n70), .A2(n71), .A3(n72), .A4(n73), .ZN(n69) );
  NOR4_X1 U10 ( .A1(n3), .A2(N59), .A3(n22), .A4(n78), .ZN(n75) );
  AOI22_X1 U11 ( .A1(n55), .A2(n100), .B1(n88), .B2(n28), .ZN(n93) );
  INV_X1 U12 ( .A(n79), .ZN(n28) );
  NAND2_X1 U13 ( .A1(n55), .A2(n99), .ZN(n72) );
  NAND2_X1 U14 ( .A1(n98), .A2(n100), .ZN(n59) );
  NOR2_X1 U15 ( .A1(n88), .A2(n72), .ZN(N21) );
  OAI211_X1 U16 ( .C1(n29), .C2(n59), .A(n93), .B(n94), .ZN(n90) );
  INV_X1 U17 ( .A(n81), .ZN(n29) );
  NAND2_X1 U18 ( .A1(n54), .A2(n80), .ZN(n92) );
  INV_X1 U19 ( .A(n52), .ZN(n25) );
  NAND2_X1 U20 ( .A1(n93), .A2(n70), .ZN(n87) );
  NAND2_X1 U21 ( .A1(n98), .A2(n99), .ZN(n77) );
  INV_X1 U22 ( .A(n71), .ZN(n21) );
  INV_X1 U23 ( .A(n54), .ZN(n22) );
  INV_X1 U24 ( .A(n76), .ZN(n27) );
  INV_X1 U25 ( .A(n94), .ZN(n20) );
  INV_X1 U26 ( .A(n68), .ZN(n10) );
  AOI22_X1 U27 ( .A1(addr_a[0]), .A2(n62), .B1(n2), .B2(n63), .ZN(n68) );
  NOR2_X1 U28 ( .A1(n77), .A2(reset), .ZN(wr_en_a) );
  NOR2_X1 U29 ( .A1(n39), .A2(state[3]), .ZN(n55) );
  NOR4_X1 U30 ( .A1(start), .A2(loadVector), .A3(loadMatrix), .A4(n80), .ZN(
        n83) );
  OAI222_X1 U31 ( .A1(n81), .A2(n24), .B1(reset), .B2(n82), .C1(N66), .C2(n19), 
        .ZN(N20) );
  INV_X1 U32 ( .A(wr_en_x), .ZN(n24) );
  NOR3_X1 U33 ( .A1(n83), .A2(n3), .A3(n21), .ZN(n82) );
  INV_X1 U34 ( .A(wr_en_a), .ZN(n19) );
  OAI21_X1 U35 ( .B1(state[1]), .B2(state[0]), .A(n55), .ZN(n52) );
  OAI22_X1 U36 ( .A1(addr_y[0]), .A2(n52), .B1(n25), .B2(n22), .ZN(n50) );
  AOI22_X1 U37 ( .A1(n81), .A2(n27), .B1(n92), .B2(start), .ZN(n94) );
  NOR2_X1 U38 ( .A1(state[3]), .A2(state[2]), .ZN(n98) );
  OAI22_X1 U39 ( .A1(loadVector), .A2(n80), .B1(n8), .B2(n72), .ZN(n97) );
  INV_X1 U40 ( .A(n88), .ZN(n8) );
  NOR2_X1 U41 ( .A1(n41), .A2(state[1]), .ZN(n99) );
  NOR2_X1 U42 ( .A1(n72), .A2(reset), .ZN(wr_en_y) );
  NOR2_X1 U43 ( .A1(n40), .A2(state[0]), .ZN(n100) );
  NOR2_X1 U44 ( .A1(n59), .A2(reset), .ZN(wr_en_x) );
  OAI21_X1 U45 ( .B1(n48), .B2(n44), .A(n49), .ZN(N56) );
  NAND4_X1 U46 ( .A1(addr_y[1]), .A2(addr_y[0]), .A3(n25), .A4(n44), .ZN(n49)
         );
  AOI21_X1 U47 ( .B1(n25), .B2(n46), .A(n50), .ZN(n48) );
  OAI21_X1 U48 ( .B1(addr_y[0]), .B2(n52), .A(n53), .ZN(N54) );
  AOI21_X1 U49 ( .B1(n95), .B2(n96), .A(reset), .ZN(N17) );
  AOI211_X1 U50 ( .C1(loadMatrix), .C2(n92), .A(n97), .B(n18), .ZN(n96) );
  AOI211_X1 U51 ( .C1(n29), .C2(n23), .A(n20), .B(n87), .ZN(n95) );
  INV_X1 U52 ( .A(n77), .ZN(n18) );
  NAND2_X1 U53 ( .A1(state[1]), .A2(n55), .ZN(n79) );
  OAI21_X1 U54 ( .B1(n7), .B2(n46), .A(n51), .ZN(N55) );
  INV_X1 U55 ( .A(n50), .ZN(n7) );
  OAI21_X1 U56 ( .B1(n17), .B2(n42), .A(n56), .ZN(N46) );
  NOR2_X1 U57 ( .A1(addr_x[0]), .A2(n17), .ZN(N44) );
  AOI21_X1 U58 ( .B1(n39), .B2(n4), .A(n5), .ZN(n3) );
  XNOR2_X1 U59 ( .A(n41), .B(state[1]), .ZN(n4) );
  NOR2_X1 U60 ( .A1(n17), .A2(n58), .ZN(N45) );
  XNOR2_X1 U61 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n58) );
  NOR2_X1 U62 ( .A1(reset), .A2(n86), .ZN(N19) );
  NOR3_X1 U63 ( .A1(n87), .A2(N21), .A3(n26), .ZN(n86) );
  INV_X1 U64 ( .A(n73), .ZN(n26) );
  NOR2_X1 U65 ( .A1(reset), .A2(n89), .ZN(N18) );
  NOR4_X1 U66 ( .A1(n90), .A2(n91), .A3(n9), .A4(n21), .ZN(n89) );
  INV_X1 U67 ( .A(n72), .ZN(n9) );
  AND3_X1 U68 ( .A1(loadVector), .A2(n30), .A3(n92), .ZN(n91) );
  INV_X1 U69 ( .A(n61), .ZN(n15) );
  AOI22_X1 U70 ( .A1(addr_a[5]), .A2(n62), .B1(N30), .B2(n63), .ZN(n61) );
  INV_X1 U71 ( .A(n66), .ZN(n12) );
  AOI22_X1 U72 ( .A1(addr_a[2]), .A2(n62), .B1(N27), .B2(n63), .ZN(n66) );
  INV_X1 U73 ( .A(n67), .ZN(n11) );
  AOI22_X1 U74 ( .A1(addr_a[1]), .A2(n62), .B1(N26), .B2(n63), .ZN(n67) );
  INV_X1 U75 ( .A(n65), .ZN(n13) );
  AOI22_X1 U76 ( .A1(addr_a[3]), .A2(n62), .B1(N28), .B2(n63), .ZN(n65) );
  INV_X1 U77 ( .A(n64), .ZN(n14) );
  AOI22_X1 U78 ( .A1(addr_a[4]), .A2(n62), .B1(N29), .B2(n63), .ZN(n64) );
  INV_X1 U79 ( .A(loadMatrix), .ZN(n30) );
  XOR2_X1 U80 ( .A(\add_103/carry[5] ), .B(addr_a[5]), .Z(N30) );
  AND3_X1 U81 ( .A1(addr_a[1]), .A2(addr_a[0]), .A3(addr_a[2]), .ZN(n6) );
  NAND4_X1 U90 ( .A1(addr_a[4]), .A2(addr_a[3]), .A3(addr_a[5]), .A4(n6), .ZN(
        N66) );
endmodule


module mvm_8_1_8_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a, wr_en_y, clear_acc;
  wire   [2:0] addr_x;
  wire   [5:0] addr_a;
  wire   [2:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a(addr_a), .wr_en_a(wr_en_a), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .clear_acc(clear_acc), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a(addr_a), .wr_en_a(wr_en_a), .clear_acc(
        clear_acc), .addr_y(addr_y), .wr_en_y(wr_en_y), .done(done), 
        .loadMatrix(loadMatrix), .loadVector(loadVector) );
endmodule

