include "s_thakkar_mvm_16_16_8_1.sv";
// Testbench, with parameters k=16, p=16, b=8, g=1

//This Test bench shows values on normal computation and in the next cycle only the vector is updated keeping the matrix same
 module tb1();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1;data_in = 65;
@(posedge clk);
#1;data_in = 66;
@(posedge clk);
#1;data_in = 67;
@(posedge clk);
#1;data_in = 68;
@(posedge clk);
#1;data_in = 69;
@(posedge clk);
#1;data_in = 70;
@(posedge clk);
#1;data_in = 71;
@(posedge clk);
#1;data_in = 72;
@(posedge clk);
#1;data_in = 73;
@(posedge clk);
#1;data_in = 74;
@(posedge clk);
#1;data_in = 75;
@(posedge clk);
#1;data_in = 76;
@(posedge clk);
#1;data_in = 77;
@(posedge clk);
#1;data_in = 78;
@(posedge clk);
#1;data_in = 79;
@(posedge clk);
#1;data_in = 80;
@(posedge clk);
#1;data_in = 81;
@(posedge clk);
#1;data_in = 82;
@(posedge clk);
#1;data_in = 83;
@(posedge clk);
#1;data_in = 84;
@(posedge clk);
#1;data_in = 85;
@(posedge clk);
#1;data_in = 86;
@(posedge clk);
#1;data_in = 87;
@(posedge clk);
#1;data_in = 88;
@(posedge clk);
#1;data_in = 89;
@(posedge clk);
#1;data_in = 90;
@(posedge clk);
#1;data_in = 91;
@(posedge clk);
#1;data_in = 92;
@(posedge clk);
#1;data_in = 93;
@(posedge clk);
#1;data_in = 94;
@(posedge clk);
#1;data_in = 95;
@(posedge clk);
#1;data_in = 96;
@(posedge clk);
#1;data_in = 97;
@(posedge clk);
#1;data_in = 98;
@(posedge clk);
#1;data_in = 99;
@(posedge clk);
#1;data_in = 100;
@(posedge clk);
#1;data_in = 101;
@(posedge clk);
#1;data_in = 102;
@(posedge clk);
#1;data_in = 103;
@(posedge clk);
#1;data_in = 104;
@(posedge clk);
#1;data_in = 105;
@(posedge clk);
#1;data_in = 106;
@(posedge clk);
#1;data_in = 107;
@(posedge clk);
#1;data_in = 108;
@(posedge clk);
#1;data_in = 109;
@(posedge clk);
#1;data_in = 110;
@(posedge clk);
#1;data_in = 111;
@(posedge clk);
#1;data_in = 112;
@(posedge clk);
#1;data_in = 113;
@(posedge clk);
#1;data_in = 114;
@(posedge clk);
#1;data_in = 115;
@(posedge clk);
#1;data_in = 116;
@(posedge clk);
#1;data_in = 117;
@(posedge clk);
#1;data_in = 118;
@(posedge clk);
#1;data_in = 119;
@(posedge clk);
#1;data_in = 120;
@(posedge clk);
#1;data_in = 121;
@(posedge clk);
#1;data_in = 122;
@(posedge clk);
#1;data_in = 123;
@(posedge clk);
#1;data_in = 124;
@(posedge clk);
#1;data_in = 125;
@(posedge clk);
#1;data_in = 126;
@(posedge clk);
#1;data_in = 127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1;data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1;data_in = 65;
@(posedge clk);
#1;data_in = 66;
@(posedge clk);
#1;data_in = 67;
@(posedge clk);
#1;data_in = 68;
@(posedge clk);
#1;data_in = 69;
@(posedge clk);
#1;data_in = 70;
@(posedge clk);
#1;data_in = 71;
@(posedge clk);
#1;data_in = 72;
@(posedge clk);
#1;data_in = 73;
@(posedge clk);
#1;data_in = 74;
@(posedge clk);
#1;data_in = 75;
@(posedge clk);
#1;data_in = 76;
@(posedge clk);
#1;data_in = 77;
@(posedge clk);
#1;data_in = 78;
@(posedge clk);
#1;data_in = 79;
@(posedge clk);
#1;data_in = 80;
@(posedge clk);
#1;data_in = 81;
@(posedge clk);
#1;data_in = 82;
@(posedge clk);
#1;data_in = 83;
@(posedge clk);
#1;data_in = 84;
@(posedge clk);
#1;data_in = 85;
@(posedge clk);
#1;data_in = 86;
@(posedge clk);
#1;data_in = 87;
@(posedge clk);
#1;data_in = 88;
@(posedge clk);
#1;data_in = 89;
@(posedge clk);
#1;data_in = 90;
@(posedge clk);
#1;data_in = 91;
@(posedge clk);
#1;data_in = 92;
@(posedge clk);
#1;data_in = 93;
@(posedge clk);
#1;data_in = 94;
@(posedge clk);
#1;data_in = 95;
@(posedge clk);
#1;data_in = 96;
@(posedge clk);
#1;data_in = 97;
@(posedge clk);
#1;data_in = 98;
@(posedge clk);
#1;data_in = 99;
@(posedge clk);
#1;data_in = 100;
@(posedge clk);
#1;data_in = 101;
@(posedge clk);
#1;data_in = 102;
@(posedge clk);
#1;data_in = 103;
@(posedge clk);
#1;data_in = 104;
@(posedge clk);
#1;data_in = 105;
@(posedge clk);
#1;data_in = 106;
@(posedge clk);
#1;data_in = 107;
@(posedge clk);
#1;data_in = 108;
@(posedge clk);
#1;data_in = 109;
@(posedge clk);
#1;data_in = 110;
@(posedge clk);
#1;data_in = 111;
@(posedge clk);
#1;data_in = 112;
@(posedge clk);
#1;data_in = 113;
@(posedge clk);
#1;data_in = 114;
@(posedge clk);
#1;data_in = 115;
@(posedge clk);
#1;data_in = 116;
@(posedge clk);
#1;data_in = 117;
@(posedge clk);
#1;data_in = 118;
@(posedge clk);
#1;data_in = 119;
@(posedge clk);
#1;data_in = 120;
@(posedge clk);
#1;data_in = 121;
@(posedge clk);
#1;data_in = 122;
@(posedge clk);
#1;data_in = 123;
@(posedge clk);
#1;data_in = 124;
@(posedge clk);
#1;data_in = 125;
@(posedge clk);
#1;data_in = 126;
@(posedge clk);
#1;data_in = 127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb1");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadVector=1;
@(posedge clk);
#1; loadVector=0;
data_in = 1;
@(posedge clk);
#1;data_in = -3;
@(posedge clk);
#1;data_in = -4;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
#1;data_in = -10;
@(posedge clk);
#1;data_in = -11;
@(posedge clk);
#1;data_in = -12;
@(posedge clk);
#1;data_in = -13;
@(posedge clk);
#1;data_in = -14;
@(posedge clk);
#1;data_in = -15;
@(posedge clk);
#1;data_in = -16;
@(posedge clk);
#1;data_in = -17;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
//This testbench incorporates two iterations in the first iteration the values are computed according to the values and in the next iteration only the Matrix is updated keeping vector
module tb2();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start = 0; reset = 1;data_in=8'bx;
@(posedge clk);
#1; reset=0;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge clk);
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1;data_in = 65;
@(posedge clk);
#1;data_in = 66;
@(posedge clk);
#1;data_in = 67;
@(posedge clk);
#1;data_in = 68;
@(posedge clk);
#1;data_in = 69;
@(posedge clk);
#1;data_in = 70;
@(posedge clk);
#1;data_in = 71;
@(posedge clk);
#1;data_in = 72;
@(posedge clk);
#1;data_in = 73;
@(posedge clk);
#1;data_in = 74;
@(posedge clk);
#1;data_in = 75;
@(posedge clk);
#1;data_in = 76;
@(posedge clk);
#1;data_in = 77;
@(posedge clk);
#1;data_in = 78;
@(posedge clk);
#1;data_in = 79;
@(posedge clk);
#1;data_in = 80;
@(posedge clk);
#1;data_in = 81;
@(posedge clk);
#1;data_in = 82;
@(posedge clk);
#1;data_in = 83;
@(posedge clk);
#1;data_in = 84;
@(posedge clk);
#1;data_in = 85;
@(posedge clk);
#1;data_in = 86;
@(posedge clk);
#1;data_in = 87;
@(posedge clk);
#1;data_in = 88;
@(posedge clk);
#1;data_in = 89;
@(posedge clk);
#1;data_in = 90;
@(posedge clk);
#1;data_in = 91;
@(posedge clk);
#1;data_in = 92;
@(posedge clk);
#1;data_in = 93;
@(posedge clk);
#1;data_in = 94;
@(posedge clk);
#1;data_in = 95;
@(posedge clk);
#1;data_in = 96;
@(posedge clk);
#1;data_in = 97;
@(posedge clk);
#1;data_in = 98;
@(posedge clk);
#1;data_in = 99;
@(posedge clk);
#1;data_in = 100;
@(posedge clk);
#1;data_in = 101;
@(posedge clk);
#1;data_in = 102;
@(posedge clk);
#1;data_in = 103;
@(posedge clk);
#1;data_in = 104;
@(posedge clk);
#1;data_in = 105;
@(posedge clk);
#1;data_in = 106;
@(posedge clk);
#1;data_in = 107;
@(posedge clk);
#1;data_in = 108;
@(posedge clk);
#1;data_in = 109;
@(posedge clk);
#1;data_in = 110;
@(posedge clk);
#1;data_in = 111;
@(posedge clk);
#1;data_in = 112;
@(posedge clk);
#1;data_in = 113;
@(posedge clk);
#1;data_in = 114;
@(posedge clk);
#1;data_in = 115;
@(posedge clk);
#1;data_in = 116;
@(posedge clk);
#1;data_in = 117;
@(posedge clk);
#1;data_in = 118;
@(posedge clk);
#1;data_in = 119;
@(posedge clk);
#1;data_in = 120;
@(posedge clk);
#1;data_in = 121;
@(posedge clk);
#1;data_in = 122;
@(posedge clk);
#1;data_in = 123;
@(posedge clk);
#1;data_in = 124;
@(posedge clk);
#1;data_in = 125;
@(posedge clk);
#1;data_in = 126;
@(posedge clk);
#1;data_in = 127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1;data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1;data_in = 65;
@(posedge clk);
#1;data_in = 66;
@(posedge clk);
#1;data_in = 67;
@(posedge clk);
#1;data_in = 68;
@(posedge clk);
#1;data_in = 69;
@(posedge clk);
#1;data_in = 70;
@(posedge clk);
#1;data_in = 71;
@(posedge clk);
#1;data_in = 72;
@(posedge clk);
#1;data_in = 73;
@(posedge clk);
#1;data_in = 74;
@(posedge clk);
#1;data_in = 75;
@(posedge clk);
#1;data_in = 76;
@(posedge clk);
#1;data_in = 77;
@(posedge clk);
#1;data_in = 78;
@(posedge clk);
#1;data_in = 79;
@(posedge clk);
#1;data_in = 80;
@(posedge clk);
#1;data_in = 81;
@(posedge clk);
#1;data_in = 82;
@(posedge clk);
#1;data_in = 83;
@(posedge clk);
#1;data_in = 84;
@(posedge clk);
#1;data_in = 85;
@(posedge clk);
#1;data_in = 86;
@(posedge clk);
#1;data_in = 87;
@(posedge clk);
#1;data_in = 88;
@(posedge clk);
#1;data_in = 89;
@(posedge clk);
#1;data_in = 90;
@(posedge clk);
#1;data_in = 91;
@(posedge clk);
#1;data_in = 92;
@(posedge clk);
#1;data_in = 93;
@(posedge clk);
#1;data_in = 94;
@(posedge clk);
#1;data_in = 95;
@(posedge clk);
#1;data_in = 96;
@(posedge clk);
#1;data_in = 97;
@(posedge clk);
#1;data_in = 98;
@(posedge clk);
#1;data_in = 99;
@(posedge clk);
#1;data_in = 100;
@(posedge clk);
#1;data_in = 101;
@(posedge clk);
#1;data_in = 102;
@(posedge clk);
#1;data_in = 103;
@(posedge clk);
#1;data_in = 104;
@(posedge clk);
#1;data_in = 105;
@(posedge clk);
#1;data_in = 106;
@(posedge clk);
#1;data_in = 107;
@(posedge clk);
#1;data_in = 108;
@(posedge clk);
#1;data_in = 109;
@(posedge clk);
#1;data_in = 110;
@(posedge clk);
#1;data_in = 111;
@(posedge clk);
#1;data_in = 112;
@(posedge clk);
#1;data_in = 113;
@(posedge clk);
#1;data_in = 114;
@(posedge clk);
#1;data_in = 115;
@(posedge clk);
#1;data_in = 116;
@(posedge clk);
#1;data_in = 117;
@(posedge clk);
#1;data_in = 118;
@(posedge clk);
#1;data_in = 119;
@(posedge clk);
#1;data_in = 120;
@(posedge clk);
#1;data_in = 121;
@(posedge clk);
#1;data_in = 122;
@(posedge clk);
#1;data_in = 123;
@(posedge clk);
#1;data_in = 124;
@(posedge clk);
#1;data_in = 125;
@(posedge clk);
#1;data_in = 126;
@(posedge clk);
#1;data_in = 127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb2");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0;
data_in = 1;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
#1;data_in = -10;
@(posedge clk);
#1;data_in = -11;
@(posedge clk);
#1;data_in = -12;
@(posedge clk);
#1;data_in = -13;
@(posedge clk);
#1;data_in = -14;
@(posedge clk);
#1;data_in = -15;
@(posedge clk);
#1;data_in = -16;
@(posedge clk);
#1;data_in = -17;
@(posedge clk);
#1;data_in = -18;
@(posedge clk);
#1;data_in = -19;
@(posedge clk);
#1;data_in = -20;
@(posedge clk);
#1;data_in = -21;
@(posedge clk);
#1;data_in = -22;
@(posedge clk);
#1;data_in = -23;
@(posedge clk);
#1;data_in = -24;
@(posedge clk);
#1;data_in = -25;
@(posedge clk);
#1;data_in = -26;
@(posedge clk);
#1;data_in = -27;
@(posedge clk);
#1;data_in = -28;
@(posedge clk);
#1;data_in = -29;
@(posedge clk);
#1;data_in = -30;
@(posedge clk);
#1;data_in = -31;
@(posedge clk);
#1;data_in = -32;
@(posedge clk);
#1;data_in = -33;
@(posedge clk);
#1;data_in = -34;
@(posedge clk);
#1;data_in = -35;
@(posedge clk);
#1;data_in = -36;
@(posedge clk);
#1;data_in = -37;
@(posedge clk);
#1;data_in = -38;
@(posedge clk);
#1;data_in = -39;
@(posedge clk);
#1;data_in = -40;
@(posedge clk);
#1;data_in = -41;
@(posedge clk);
#1;data_in = -42;
@(posedge clk);
#1;data_in = -43;
@(posedge clk);
#1;data_in = -44;
@(posedge clk);
#1;data_in = -45;
@(posedge clk);
#1;data_in = -46;
@(posedge clk);
#1;data_in = -47;
@(posedge clk);
#1;data_in = -48;
@(posedge clk);
#1;data_in = -49;
@(posedge clk);
#1;data_in = -50;
@(posedge clk);
#1;data_in = -51;
@(posedge clk);
#1;data_in = -52;
@(posedge clk);
#1;data_in = -53;
@(posedge clk);
#1;data_in = -54;
@(posedge clk);
#1;data_in = -55;
@(posedge clk);
#1;data_in = -56;
@(posedge clk);
#1;data_in = -57;
@(posedge clk);
#1;data_in = -58;
@(posedge clk);
#1;data_in = -59;
@(posedge clk);
#1;data_in = -60;
@(posedge clk);
#1;data_in = -61;
@(posedge clk);
#1;data_in = -62;
@(posedge clk);
#1;data_in = -63;
@(posedge clk);
#1;data_in = -64;
@(posedge clk);
#1;data_in = -65;
@(posedge clk);
#1;data_in = -66;
@(posedge clk);
#1;data_in = -67;
@(posedge clk);
#1;data_in = -68;
@(posedge clk);
#1;data_in = -69;
@(posedge clk);
#1;data_in = -70;
@(posedge clk);
#1;data_in = -71;
@(posedge clk);
#1;data_in = -72;
@(posedge clk);
#1;data_in = -73;
@(posedge clk);
#1;data_in = -74;
@(posedge clk);
#1;data_in = -75;
@(posedge clk);
#1;data_in = -76;
@(posedge clk);
#1;data_in = -77;
@(posedge clk);
#1;data_in = -78;
@(posedge clk);
#1;data_in = -79;
@(posedge clk);
#1;data_in = -80;
@(posedge clk);
#1;data_in = -81;
@(posedge clk);
#1;data_in = -82;
@(posedge clk);
#1;data_in = -83;
@(posedge clk);
#1;data_in = -84;
@(posedge clk);
#1;data_in = -85;
@(posedge clk);
#1;data_in = -86;
@(posedge clk);
#1;data_in = -87;
@(posedge clk);
#1;data_in = -88;
@(posedge clk);
#1;data_in = -89;
@(posedge clk);
#1;data_in = -90;
@(posedge clk);
#1;data_in = -91;
@(posedge clk);
#1;data_in = -92;
@(posedge clk);
#1;data_in = -93;
@(posedge clk);
#1;data_in = -94;
@(posedge clk);
#1;data_in = -95;
@(posedge clk);
#1;data_in = -96;
@(posedge clk);
#1;data_in = -97;
@(posedge clk);
#1;data_in = -98;
@(posedge clk);
#1;data_in = -99;
@(posedge clk);
#1;data_in = -100;
@(posedge clk);
#1;data_in = -101;
@(posedge clk);
#1;data_in = -102;
@(posedge clk);
#1;data_in = -103;
@(posedge clk);
#1;data_in = -104;
@(posedge clk);
#1;data_in = -105;
@(posedge clk);
#1;data_in = -106;
@(posedge clk);
#1;data_in = -107;
@(posedge clk);
#1;data_in = -108;
@(posedge clk);
#1;data_in = -109;
@(posedge clk);
#1;data_in = -110;
@(posedge clk);
#1;data_in = -111;
@(posedge clk);
#1;data_in = -112;
@(posedge clk);
#1;data_in = -113;
@(posedge clk);
#1;data_in = -114;
@(posedge clk);
#1;data_in = -115;
@(posedge clk);
#1;data_in = -116;
@(posedge clk);
#1;data_in = -117;
@(posedge clk);
#1;data_in = -118;
@(posedge clk);
#1;data_in = -119;
@(posedge clk);
#1;data_in = -120;
@(posedge clk);
#1;data_in = -121;
@(posedge clk);
#1;data_in = -122;
@(posedge clk);
#1;data_in = -123;
@(posedge clk);
#1;data_in = -124;
@(posedge clk);
#1;data_in = -125;
@(posedge clk);
#1;data_in = -126;
@(posedge clk);
#1;data_in = -127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1;data_in = -1;
@(posedge clk);
#1;data_in = -2;
@(posedge clk);
#1;data_in = -3;
@(posedge clk);
#1;data_in = -4;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
#1;data_in = -10;
@(posedge clk);
#1;data_in = -11;
@(posedge clk);
#1;data_in = -12;
@(posedge clk);
#1;data_in = -13;
@(posedge clk);
#1;data_in = -14;
@(posedge clk);
#1;data_in = -15;
@(posedge clk);
#1;data_in = -16;
@(posedge clk);
#1;data_in = -17;
@(posedge clk);
#1;data_in = -18;
@(posedge clk);
#1;data_in = -19;
@(posedge clk);
#1;data_in = -20;
@(posedge clk);
#1;data_in = -21;
@(posedge clk);
#1;data_in = -22;
@(posedge clk);
#1;data_in = -23;
@(posedge clk);
#1;data_in = -24;
@(posedge clk);
#1;data_in = -25;
@(posedge clk);
#1;data_in = -26;
@(posedge clk);
#1;data_in = -27;
@(posedge clk);
#1;data_in = -28;
@(posedge clk);
#1;data_in = -29;
@(posedge clk);
#1;data_in = -30;
@(posedge clk);
#1;data_in = -31;
@(posedge clk);
#1;data_in = -32;
@(posedge clk);
#1;data_in = -33;
@(posedge clk);
#1;data_in = -34;
@(posedge clk);
#1;data_in = -35;
@(posedge clk);
#1;data_in = -36;
@(posedge clk);
#1;data_in = -37;
@(posedge clk);
#1;data_in = -38;
@(posedge clk);
#1;data_in = -39;
@(posedge clk);
#1;data_in = -40;
@(posedge clk);
#1;data_in = -41;
@(posedge clk);
#1;data_in = -42;
@(posedge clk);
#1;data_in = -43;
@(posedge clk);
#1;data_in = -44;
@(posedge clk);
#1;data_in = -45;
@(posedge clk);
#1;data_in = -46;
@(posedge clk);
#1;data_in = -47;
@(posedge clk);
#1;data_in = -48;
@(posedge clk);
#1;data_in = -49;
@(posedge clk);
#1;data_in = -50;
@(posedge clk);
#1;data_in = -51;
@(posedge clk);
#1;data_in = -52;
@(posedge clk);
#1;data_in = -53;
@(posedge clk);
#1;data_in = -54;
@(posedge clk);
#1;data_in = -55;
@(posedge clk);
#1;data_in = -56;
@(posedge clk);
#1;data_in = -57;
@(posedge clk);
#1;data_in = -58;
@(posedge clk);
#1;data_in = -59;
@(posedge clk);
#1;data_in = -60;
@(posedge clk);
#1;data_in = -61;
@(posedge clk);
#1;data_in = -62;
@(posedge clk);
#1;data_in = -63;
@(posedge clk);
#1;data_in = -64;
@(posedge clk);
#1;data_in = -65;
@(posedge clk);
#1;data_in = -66;
@(posedge clk);
#1;data_in = -67;
@(posedge clk);
#1;data_in = -68;
@(posedge clk);
#1;data_in = -69;
@(posedge clk);
#1;data_in = -70;
@(posedge clk);
#1;data_in = -71;
@(posedge clk);
#1;data_in = -72;
@(posedge clk);
#1;data_in = -73;
@(posedge clk);
#1;data_in = -74;
@(posedge clk);
#1;data_in = -75;
@(posedge clk);
#1;data_in = -76;
@(posedge clk);
#1;data_in = -77;
@(posedge clk);
#1;data_in = -78;
@(posedge clk);
#1;data_in = -79;
@(posedge clk);
#1;data_in = -80;
@(posedge clk);
#1;data_in = -81;
@(posedge clk);
#1;data_in = -82;
@(posedge clk);
#1;data_in = -83;
@(posedge clk);
#1;data_in = -84;
@(posedge clk);
#1;data_in = -85;
@(posedge clk);
#1;data_in = -86;
@(posedge clk);
#1;data_in = -87;
@(posedge clk);
#1;data_in = -88;
@(posedge clk);
#1;data_in = -89;
@(posedge clk);
#1;data_in = -90;
@(posedge clk);
#1;data_in = -91;
@(posedge clk);
#1;data_in = -92;
@(posedge clk);
#1;data_in = -93;
@(posedge clk);
#1;data_in = -94;
@(posedge clk);
#1;data_in = -95;
@(posedge clk);
#1;data_in = -96;
@(posedge clk);
#1;data_in = -97;
@(posedge clk);
#1;data_in = -98;
@(posedge clk);
#1;data_in = -99;
@(posedge clk);
#1;data_in = -100;
@(posedge clk);
#1;data_in = -101;
@(posedge clk);
#1;data_in = -102;
@(posedge clk);
#1;data_in = -103;
@(posedge clk);
#1;data_in = -104;
@(posedge clk);
#1;data_in = -105;
@(posedge clk);
#1;data_in = -106;
@(posedge clk);
#1;data_in = -107;
@(posedge clk);
#1;data_in = -108;
@(posedge clk);
#1;data_in = -109;
@(posedge clk);
#1;data_in = -110;
@(posedge clk);
#1;data_in = -111;
@(posedge clk);
#1;data_in = -112;
@(posedge clk);
#1;data_in = -113;
@(posedge clk);
#1;data_in = -114;
@(posedge clk);
#1;data_in = -115;
@(posedge clk);
#1;data_in = -116;
@(posedge clk);
#1;data_in = -117;
@(posedge clk);
#1;data_in = -118;
@(posedge clk);
#1;data_in = -119;
@(posedge clk);
#1;data_in = -120;
@(posedge clk);
#1;data_in = -121;
@(posedge clk);
#1;data_in = -122;
@(posedge clk);
#1;data_in = -123;
@(posedge clk);
#1;data_in = -124;
@(posedge clk);
#1;data_in = -125;
@(posedge clk);
#1;data_in = -126;
@(posedge clk);
#1;data_in = -127;
@(posedge clk);
#1;data_in = 0;
@(posedge clk);
#1;data_in = -1;
@(posedge clk);
#1;data_in = -2;
@(posedge clk);
#1;data_in = -3;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=16, p=16, b=8, g=1

module tb3();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData3[271:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb3", testData3);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb3");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData3[0];
@(posedge clk);
#1;data_in = testData3[1];
@(posedge clk);
#1;data_in = testData3[2];
@(posedge clk);
#1;data_in = testData3[3];
@(posedge clk);
#1;data_in = testData3[4];
@(posedge clk);
#1;data_in = testData3[5];
@(posedge clk);
#1;data_in = testData3[6];
@(posedge clk);
#1;data_in = testData3[7];
@(posedge clk);
#1;data_in = testData3[8];
@(posedge clk);
#1;data_in = testData3[9];
@(posedge clk);
#1;data_in = testData3[10];
@(posedge clk);
#1;data_in = testData3[11];
@(posedge clk);
#1;data_in = testData3[12];
@(posedge clk);
#1;data_in = testData3[13];
@(posedge clk);
#1;data_in = testData3[14];
@(posedge clk);
#1;data_in = testData3[15];
@(posedge clk);
#1;data_in = testData3[16];
@(posedge clk);
#1;data_in = testData3[17];
@(posedge clk);
#1;data_in = testData3[18];
@(posedge clk);
#1;data_in = testData3[19];
@(posedge clk);
#1;data_in = testData3[20];
@(posedge clk);
#1;data_in = testData3[21];
@(posedge clk);
#1;data_in = testData3[22];
@(posedge clk);
#1;data_in = testData3[23];
@(posedge clk);
#1;data_in = testData3[24];
@(posedge clk);
#1;data_in = testData3[25];
@(posedge clk);
#1;data_in = testData3[26];
@(posedge clk);
#1;data_in = testData3[27];
@(posedge clk);
#1;data_in = testData3[28];
@(posedge clk);
#1;data_in = testData3[29];
@(posedge clk);
#1;data_in = testData3[30];
@(posedge clk);
#1;data_in = testData3[31];
@(posedge clk);
#1;data_in = testData3[32];
@(posedge clk);
#1;data_in = testData3[33];
@(posedge clk);
#1;data_in = testData3[34];
@(posedge clk);
#1;data_in = testData3[35];
@(posedge clk);
#1;data_in = testData3[36];
@(posedge clk);
#1;data_in = testData3[37];
@(posedge clk);
#1;data_in = testData3[38];
@(posedge clk);
#1;data_in = testData3[39];
@(posedge clk);
#1;data_in = testData3[40];
@(posedge clk);
#1;data_in = testData3[41];
@(posedge clk);
#1;data_in = testData3[42];
@(posedge clk);
#1;data_in = testData3[43];
@(posedge clk);
#1;data_in = testData3[44];
@(posedge clk);
#1;data_in = testData3[45];
@(posedge clk);
#1;data_in = testData3[46];
@(posedge clk);
#1;data_in = testData3[47];
@(posedge clk);
#1;data_in = testData3[48];
@(posedge clk);
#1;data_in = testData3[49];
@(posedge clk);
#1;data_in = testData3[50];
@(posedge clk);
#1;data_in = testData3[51];
@(posedge clk);
#1;data_in = testData3[52];
@(posedge clk);
#1;data_in = testData3[53];
@(posedge clk);
#1;data_in = testData3[54];
@(posedge clk);
#1;data_in = testData3[55];
@(posedge clk);
#1;data_in = testData3[56];
@(posedge clk);
#1;data_in = testData3[57];
@(posedge clk);
#1;data_in = testData3[58];
@(posedge clk);
#1;data_in = testData3[59];
@(posedge clk);
#1;data_in = testData3[60];
@(posedge clk);
#1;data_in = testData3[61];
@(posedge clk);
#1;data_in = testData3[62];
@(posedge clk);
#1;data_in = testData3[63];
@(posedge clk);
#1;data_in = testData3[64];
@(posedge clk);
#1;data_in = testData3[65];
@(posedge clk);
#1;data_in = testData3[66];
@(posedge clk);
#1;data_in = testData3[67];
@(posedge clk);
#1;data_in = testData3[68];
@(posedge clk);
#1;data_in = testData3[69];
@(posedge clk);
#1;data_in = testData3[70];
@(posedge clk);
#1;data_in = testData3[71];
@(posedge clk);
#1;data_in = testData3[72];
@(posedge clk);
#1;data_in = testData3[73];
@(posedge clk);
#1;data_in = testData3[74];
@(posedge clk);
#1;data_in = testData3[75];
@(posedge clk);
#1;data_in = testData3[76];
@(posedge clk);
#1;data_in = testData3[77];
@(posedge clk);
#1;data_in = testData3[78];
@(posedge clk);
#1;data_in = testData3[79];
@(posedge clk);
#1;data_in = testData3[80];
@(posedge clk);
#1;data_in = testData3[81];
@(posedge clk);
#1;data_in = testData3[82];
@(posedge clk);
#1;data_in = testData3[83];
@(posedge clk);
#1;data_in = testData3[84];
@(posedge clk);
#1;data_in = testData3[85];
@(posedge clk);
#1;data_in = testData3[86];
@(posedge clk);
#1;data_in = testData3[87];
@(posedge clk);
#1;data_in = testData3[88];
@(posedge clk);
#1;data_in = testData3[89];
@(posedge clk);
#1;data_in = testData3[90];
@(posedge clk);
#1;data_in = testData3[91];
@(posedge clk);
#1;data_in = testData3[92];
@(posedge clk);
#1;data_in = testData3[93];
@(posedge clk);
#1;data_in = testData3[94];
@(posedge clk);
#1;data_in = testData3[95];
@(posedge clk);
#1;data_in = testData3[96];
@(posedge clk);
#1;data_in = testData3[97];
@(posedge clk);
#1;data_in = testData3[98];
@(posedge clk);
#1;data_in = testData3[99];
@(posedge clk);
#1;data_in = testData3[100];
@(posedge clk);
#1;data_in = testData3[101];
@(posedge clk);
#1;data_in = testData3[102];
@(posedge clk);
#1;data_in = testData3[103];
@(posedge clk);
#1;data_in = testData3[104];
@(posedge clk);
#1;data_in = testData3[105];
@(posedge clk);
#1;data_in = testData3[106];
@(posedge clk);
#1;data_in = testData3[107];
@(posedge clk);
#1;data_in = testData3[108];
@(posedge clk);
#1;data_in = testData3[109];
@(posedge clk);
#1;data_in = testData3[110];
@(posedge clk);
#1;data_in = testData3[111];
@(posedge clk);
#1;data_in = testData3[112];
@(posedge clk);
#1;data_in = testData3[113];
@(posedge clk);
#1;data_in = testData3[114];
@(posedge clk);
#1;data_in = testData3[115];
@(posedge clk);
#1;data_in = testData3[116];
@(posedge clk);
#1;data_in = testData3[117];
@(posedge clk);
#1;data_in = testData3[118];
@(posedge clk);
#1;data_in = testData3[119];
@(posedge clk);
#1;data_in = testData3[120];
@(posedge clk);
#1;data_in = testData3[121];
@(posedge clk);
#1;data_in = testData3[122];
@(posedge clk);
#1;data_in = testData3[123];
@(posedge clk);
#1;data_in = testData3[124];
@(posedge clk);
#1;data_in = testData3[125];
@(posedge clk);
#1;data_in = testData3[126];
@(posedge clk);
#1;data_in = testData3[127];
@(posedge clk);
#1;data_in = testData3[128];
@(posedge clk);
#1;data_in = testData3[129];
@(posedge clk);
#1;data_in = testData3[130];
@(posedge clk);
#1;data_in = testData3[131];
@(posedge clk);
#1;data_in = testData3[132];
@(posedge clk);
#1;data_in = testData3[133];
@(posedge clk);
#1;data_in = testData3[134];
@(posedge clk);
#1;data_in = testData3[135];
@(posedge clk);
#1;data_in = testData3[136];
@(posedge clk);
#1;data_in = testData3[137];
@(posedge clk);
#1;data_in = testData3[138];
@(posedge clk);
#1;data_in = testData3[139];
@(posedge clk);
#1;data_in = testData3[140];
@(posedge clk);
#1;data_in = testData3[141];
@(posedge clk);
#1;data_in = testData3[142];
@(posedge clk);
#1;data_in = testData3[143];
@(posedge clk);
#1;data_in = testData3[144];
@(posedge clk);
#1;data_in = testData3[145];
@(posedge clk);
#1;data_in = testData3[146];
@(posedge clk);
#1;data_in = testData3[147];
@(posedge clk);
#1;data_in = testData3[148];
@(posedge clk);
#1;data_in = testData3[149];
@(posedge clk);
#1;data_in = testData3[150];
@(posedge clk);
#1;data_in = testData3[151];
@(posedge clk);
#1;data_in = testData3[152];
@(posedge clk);
#1;data_in = testData3[153];
@(posedge clk);
#1;data_in = testData3[154];
@(posedge clk);
#1;data_in = testData3[155];
@(posedge clk);
#1;data_in = testData3[156];
@(posedge clk);
#1;data_in = testData3[157];
@(posedge clk);
#1;data_in = testData3[158];
@(posedge clk);
#1;data_in = testData3[159];
@(posedge clk);
#1;data_in = testData3[160];
@(posedge clk);
#1;data_in = testData3[161];
@(posedge clk);
#1;data_in = testData3[162];
@(posedge clk);
#1;data_in = testData3[163];
@(posedge clk);
#1;data_in = testData3[164];
@(posedge clk);
#1;data_in = testData3[165];
@(posedge clk);
#1;data_in = testData3[166];
@(posedge clk);
#1;data_in = testData3[167];
@(posedge clk);
#1;data_in = testData3[168];
@(posedge clk);
#1;data_in = testData3[169];
@(posedge clk);
#1;data_in = testData3[170];
@(posedge clk);
#1;data_in = testData3[171];
@(posedge clk);
#1;data_in = testData3[172];
@(posedge clk);
#1;data_in = testData3[173];
@(posedge clk);
#1;data_in = testData3[174];
@(posedge clk);
#1;data_in = testData3[175];
@(posedge clk);
#1;data_in = testData3[176];
@(posedge clk);
#1;data_in = testData3[177];
@(posedge clk);
#1;data_in = testData3[178];
@(posedge clk);
#1;data_in = testData3[179];
@(posedge clk);
#1;data_in = testData3[180];
@(posedge clk);
#1;data_in = testData3[181];
@(posedge clk);
#1;data_in = testData3[182];
@(posedge clk);
#1;data_in = testData3[183];
@(posedge clk);
#1;data_in = testData3[184];
@(posedge clk);
#1;data_in = testData3[185];
@(posedge clk);
#1;data_in = testData3[186];
@(posedge clk);
#1;data_in = testData3[187];
@(posedge clk);
#1;data_in = testData3[188];
@(posedge clk);
#1;data_in = testData3[189];
@(posedge clk);
#1;data_in = testData3[190];
@(posedge clk);
#1;data_in = testData3[191];
@(posedge clk);
#1;data_in = testData3[192];
@(posedge clk);
#1;data_in = testData3[193];
@(posedge clk);
#1;data_in = testData3[194];
@(posedge clk);
#1;data_in = testData3[195];
@(posedge clk);
#1;data_in = testData3[196];
@(posedge clk);
#1;data_in = testData3[197];
@(posedge clk);
#1;data_in = testData3[198];
@(posedge clk);
#1;data_in = testData3[199];
@(posedge clk);
#1;data_in = testData3[200];
@(posedge clk);
#1;data_in = testData3[201];
@(posedge clk);
#1;data_in = testData3[202];
@(posedge clk);
#1;data_in = testData3[203];
@(posedge clk);
#1;data_in = testData3[204];
@(posedge clk);
#1;data_in = testData3[205];
@(posedge clk);
#1;data_in = testData3[206];
@(posedge clk);
#1;data_in = testData3[207];
@(posedge clk);
#1;data_in = testData3[208];
@(posedge clk);
#1;data_in = testData3[209];
@(posedge clk);
#1;data_in = testData3[210];
@(posedge clk);
#1;data_in = testData3[211];
@(posedge clk);
#1;data_in = testData3[212];
@(posedge clk);
#1;data_in = testData3[213];
@(posedge clk);
#1;data_in = testData3[214];
@(posedge clk);
#1;data_in = testData3[215];
@(posedge clk);
#1;data_in = testData3[216];
@(posedge clk);
#1;data_in = testData3[217];
@(posedge clk);
#1;data_in = testData3[218];
@(posedge clk);
#1;data_in = testData3[219];
@(posedge clk);
#1;data_in = testData3[220];
@(posedge clk);
#1;data_in = testData3[221];
@(posedge clk);
#1;data_in = testData3[222];
@(posedge clk);
#1;data_in = testData3[223];
@(posedge clk);
#1;data_in = testData3[224];
@(posedge clk);
#1;data_in = testData3[225];
@(posedge clk);
#1;data_in = testData3[226];
@(posedge clk);
#1;data_in = testData3[227];
@(posedge clk);
#1;data_in = testData3[228];
@(posedge clk);
#1;data_in = testData3[229];
@(posedge clk);
#1;data_in = testData3[230];
@(posedge clk);
#1;data_in = testData3[231];
@(posedge clk);
#1;data_in = testData3[232];
@(posedge clk);
#1;data_in = testData3[233];
@(posedge clk);
#1;data_in = testData3[234];
@(posedge clk);
#1;data_in = testData3[235];
@(posedge clk);
#1;data_in = testData3[236];
@(posedge clk);
#1;data_in = testData3[237];
@(posedge clk);
#1;data_in = testData3[238];
@(posedge clk);
#1;data_in = testData3[239];
@(posedge clk);
#1;data_in = testData3[240];
@(posedge clk);
#1;data_in = testData3[241];
@(posedge clk);
#1;data_in = testData3[242];
@(posedge clk);
#1;data_in = testData3[243];
@(posedge clk);
#1;data_in = testData3[244];
@(posedge clk);
#1;data_in = testData3[245];
@(posedge clk);
#1;data_in = testData3[246];
@(posedge clk);
#1;data_in = testData3[247];
@(posedge clk);
#1;data_in = testData3[248];
@(posedge clk);
#1;data_in = testData3[249];
@(posedge clk);
#1;data_in = testData3[250];
@(posedge clk);
#1;data_in = testData3[251];
@(posedge clk);
#1;data_in = testData3[252];
@(posedge clk);
#1;data_in = testData3[253];
@(posedge clk);
#1;data_in = testData3[254];
@(posedge clk);
#1;data_in = testData3[255];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData3[256]; 
@(posedge clk);
#1;data_in = testData3[257];
@(posedge clk);
#1;data_in = testData3[258];
@(posedge clk);
#1;data_in = testData3[259];
@(posedge clk);
#1;data_in = testData3[260];
@(posedge clk);
#1;data_in = testData3[261];
@(posedge clk);
#1;data_in = testData3[262];
@(posedge clk);
#1;data_in = testData3[263];
@(posedge clk);
#1;data_in = testData3[264];
@(posedge clk);
#1;data_in = testData3[265];
@(posedge clk);
#1;data_in = testData3[266];
@(posedge clk);
#1;data_in = testData3[267];
@(posedge clk);
#1;data_in = testData3[268];
@(posedge clk);
#1;data_in = testData3[269];
@(posedge clk);
#1;data_in = testData3[270];
@(posedge clk);
#1;data_in = testData3[271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=16, p=16, b=8, g=1

module tb4();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData4[1071:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb4", testData4);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb4");
  initial begin 
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData4[0];
@(posedge clk);
#1;data_in = testData4[1];
@(posedge clk);
#1;data_in = testData4[2];
@(posedge clk);
#1;data_in = testData4[3];
@(posedge clk);
#1;data_in = testData4[4];
@(posedge clk);
#1;data_in = testData4[5];
@(posedge clk);
#1;data_in = testData4[6];
@(posedge clk);
#1;data_in = testData4[7];
@(posedge clk);
#1;data_in = testData4[8];
@(posedge clk);
#1;data_in = testData4[9];
@(posedge clk);
#1;data_in = testData4[10];
@(posedge clk);
#1;data_in = testData4[11];
@(posedge clk);
#1;data_in = testData4[12];
@(posedge clk);
#1;data_in = testData4[13];
@(posedge clk);
#1;data_in = testData4[14];
@(posedge clk);
#1;data_in = testData4[15];
@(posedge clk);
#1;data_in = testData4[16];
@(posedge clk);
#1;data_in = testData4[17];
@(posedge clk);
#1;data_in = testData4[18];
@(posedge clk);
#1;data_in = testData4[19];
@(posedge clk);
#1;data_in = testData4[20];
@(posedge clk);
#1;data_in = testData4[21];
@(posedge clk);
#1;data_in = testData4[22];
@(posedge clk);
#1;data_in = testData4[23];
@(posedge clk);
#1;data_in = testData4[24];
@(posedge clk);
#1;data_in = testData4[25];
@(posedge clk);
#1;data_in = testData4[26];
@(posedge clk);
#1;data_in = testData4[27];
@(posedge clk);
#1;data_in = testData4[28];
@(posedge clk);
#1;data_in = testData4[29];
@(posedge clk);
#1;data_in = testData4[30];
@(posedge clk);
#1;data_in = testData4[31];
@(posedge clk);
#1;data_in = testData4[32];
@(posedge clk);
#1;data_in = testData4[33];
@(posedge clk);
#1;data_in = testData4[34];
@(posedge clk);
#1;data_in = testData4[35];
@(posedge clk);
#1;data_in = testData4[36];
@(posedge clk);
#1;data_in = testData4[37];
@(posedge clk);
#1;data_in = testData4[38];
@(posedge clk);
#1;data_in = testData4[39];
@(posedge clk);
#1;data_in = testData4[40];
@(posedge clk);
#1;data_in = testData4[41];
@(posedge clk);
#1;data_in = testData4[42];
@(posedge clk);
#1;data_in = testData4[43];
@(posedge clk);
#1;data_in = testData4[44];
@(posedge clk);
#1;data_in = testData4[45];
@(posedge clk);
#1;data_in = testData4[46];
@(posedge clk);
#1;data_in = testData4[47];
@(posedge clk);
#1;data_in = testData4[48];
@(posedge clk);
#1;data_in = testData4[49];
@(posedge clk);
#1;data_in = testData4[50];
@(posedge clk);
#1;data_in = testData4[51];
@(posedge clk);
#1;data_in = testData4[52];
@(posedge clk);
#1;data_in = testData4[53];
@(posedge clk);
#1;data_in = testData4[54];
@(posedge clk);
#1;data_in = testData4[55];
@(posedge clk);
#1;data_in = testData4[56];
@(posedge clk);
#1;data_in = testData4[57];
@(posedge clk);
#1;data_in = testData4[58];
@(posedge clk);
#1;data_in = testData4[59];
@(posedge clk);
#1;data_in = testData4[60];
@(posedge clk);
#1;data_in = testData4[61];
@(posedge clk);
#1;data_in = testData4[62];
@(posedge clk);
#1;data_in = testData4[63];
@(posedge clk);
#1;data_in = testData4[64];
@(posedge clk);
#1;data_in = testData4[65];
@(posedge clk);
#1;data_in = testData4[66];
@(posedge clk);
#1;data_in = testData4[67];
@(posedge clk);
#1;data_in = testData4[68];
@(posedge clk);
#1;data_in = testData4[69];
@(posedge clk);
#1;data_in = testData4[70];
@(posedge clk);
#1;data_in = testData4[71];
@(posedge clk);
#1;data_in = testData4[72];
@(posedge clk);
#1;data_in = testData4[73];
@(posedge clk);
#1;data_in = testData4[74];
@(posedge clk);
#1;data_in = testData4[75];
@(posedge clk);
#1;data_in = testData4[76];
@(posedge clk);
#1;data_in = testData4[77];
@(posedge clk);
#1;data_in = testData4[78];
@(posedge clk);
#1;data_in = testData4[79];
@(posedge clk);
#1;data_in = testData4[80];
@(posedge clk);
#1;data_in = testData4[81];
@(posedge clk);
#1;data_in = testData4[82];
@(posedge clk);
#1;data_in = testData4[83];
@(posedge clk);
#1;data_in = testData4[84];
@(posedge clk);
#1;data_in = testData4[85];
@(posedge clk);
#1;data_in = testData4[86];
@(posedge clk);
#1;data_in = testData4[87];
@(posedge clk);
#1;data_in = testData4[88];
@(posedge clk);
#1;data_in = testData4[89];
@(posedge clk);
#1;data_in = testData4[90];
@(posedge clk);
#1;data_in = testData4[91];
@(posedge clk);
#1;data_in = testData4[92];
@(posedge clk);
#1;data_in = testData4[93];
@(posedge clk);
#1;data_in = testData4[94];
@(posedge clk);
#1;data_in = testData4[95];
@(posedge clk);
#1;data_in = testData4[96];
@(posedge clk);
#1;data_in = testData4[97];
@(posedge clk);
#1;data_in = testData4[98];
@(posedge clk);
#1;data_in = testData4[99];
@(posedge clk);
#1;data_in = testData4[100];
@(posedge clk);
#1;data_in = testData4[101];
@(posedge clk);
#1;data_in = testData4[102];
@(posedge clk);
#1;data_in = testData4[103];
@(posedge clk);
#1;data_in = testData4[104];
@(posedge clk);
#1;data_in = testData4[105];
@(posedge clk);
#1;data_in = testData4[106];
@(posedge clk);
#1;data_in = testData4[107];
@(posedge clk);
#1;data_in = testData4[108];
@(posedge clk);
#1;data_in = testData4[109];
@(posedge clk);
#1;data_in = testData4[110];
@(posedge clk);
#1;data_in = testData4[111];
@(posedge clk);
#1;data_in = testData4[112];
@(posedge clk);
#1;data_in = testData4[113];
@(posedge clk);
#1;data_in = testData4[114];
@(posedge clk);
#1;data_in = testData4[115];
@(posedge clk);
#1;data_in = testData4[116];
@(posedge clk);
#1;data_in = testData4[117];
@(posedge clk);
#1;data_in = testData4[118];
@(posedge clk);
#1;data_in = testData4[119];
@(posedge clk);
#1;data_in = testData4[120];
@(posedge clk);
#1;data_in = testData4[121];
@(posedge clk);
#1;data_in = testData4[122];
@(posedge clk);
#1;data_in = testData4[123];
@(posedge clk);
#1;data_in = testData4[124];
@(posedge clk);
#1;data_in = testData4[125];
@(posedge clk);
#1;data_in = testData4[126];
@(posedge clk);
#1;data_in = testData4[127];
@(posedge clk);
#1;data_in = testData4[128];
@(posedge clk);
#1;data_in = testData4[129];
@(posedge clk);
#1;data_in = testData4[130];
@(posedge clk);
#1;data_in = testData4[131];
@(posedge clk);
#1;data_in = testData4[132];
@(posedge clk);
#1;data_in = testData4[133];
@(posedge clk);
#1;data_in = testData4[134];
@(posedge clk);
#1;data_in = testData4[135];
@(posedge clk);
#1;data_in = testData4[136];
@(posedge clk);
#1;data_in = testData4[137];
@(posedge clk);
#1;data_in = testData4[138];
@(posedge clk);
#1;data_in = testData4[139];
@(posedge clk);
#1;data_in = testData4[140];
@(posedge clk);
#1;data_in = testData4[141];
@(posedge clk);
#1;data_in = testData4[142];
@(posedge clk);
#1;data_in = testData4[143];
@(posedge clk);
#1;data_in = testData4[144];
@(posedge clk);
#1;data_in = testData4[145];
@(posedge clk);
#1;data_in = testData4[146];
@(posedge clk);
#1;data_in = testData4[147];
@(posedge clk);
#1;data_in = testData4[148];
@(posedge clk);
#1;data_in = testData4[149];
@(posedge clk);
#1;data_in = testData4[150];
@(posedge clk);
#1;data_in = testData4[151];
@(posedge clk);
#1;data_in = testData4[152];
@(posedge clk);
#1;data_in = testData4[153];
@(posedge clk);
#1;data_in = testData4[154];
@(posedge clk);
#1;data_in = testData4[155];
@(posedge clk);
#1;data_in = testData4[156];
@(posedge clk);
#1;data_in = testData4[157];
@(posedge clk);
#1;data_in = testData4[158];
@(posedge clk);
#1;data_in = testData4[159];
@(posedge clk);
#1;data_in = testData4[160];
@(posedge clk);
#1;data_in = testData4[161];
@(posedge clk);
#1;data_in = testData4[162];
@(posedge clk);
#1;data_in = testData4[163];
@(posedge clk);
#1;data_in = testData4[164];
@(posedge clk);
#1;data_in = testData4[165];
@(posedge clk);
#1;data_in = testData4[166];
@(posedge clk);
#1;data_in = testData4[167];
@(posedge clk);
#1;data_in = testData4[168];
@(posedge clk);
#1;data_in = testData4[169];
@(posedge clk);
#1;data_in = testData4[170];
@(posedge clk);
#1;data_in = testData4[171];
@(posedge clk);
#1;data_in = testData4[172];
@(posedge clk);
#1;data_in = testData4[173];
@(posedge clk);
#1;data_in = testData4[174];
@(posedge clk);
#1;data_in = testData4[175];
@(posedge clk);
#1;data_in = testData4[176];
@(posedge clk);
#1;data_in = testData4[177];
@(posedge clk);
#1;data_in = testData4[178];
@(posedge clk);
#1;data_in = testData4[179];
@(posedge clk);
#1;data_in = testData4[180];
@(posedge clk);
#1;data_in = testData4[181];
@(posedge clk);
#1;data_in = testData4[182];
@(posedge clk);
#1;data_in = testData4[183];
@(posedge clk);
#1;data_in = testData4[184];
@(posedge clk);
#1;data_in = testData4[185];
@(posedge clk);
#1;data_in = testData4[186];
@(posedge clk);
#1;data_in = testData4[187];
@(posedge clk);
#1;data_in = testData4[188];
@(posedge clk);
#1;data_in = testData4[189];
@(posedge clk);
#1;data_in = testData4[190];
@(posedge clk);
#1;data_in = testData4[191];
@(posedge clk);
#1;data_in = testData4[192];
@(posedge clk);
#1;data_in = testData4[193];
@(posedge clk);
#1;data_in = testData4[194];
@(posedge clk);
#1;data_in = testData4[195];
@(posedge clk);
#1;data_in = testData4[196];
@(posedge clk);
#1;data_in = testData4[197];
@(posedge clk);
#1;data_in = testData4[198];
@(posedge clk);
#1;data_in = testData4[199];
@(posedge clk);
#1;data_in = testData4[200];
@(posedge clk);
#1;data_in = testData4[201];
@(posedge clk);
#1;data_in = testData4[202];
@(posedge clk);
#1;data_in = testData4[203];
@(posedge clk);
#1;data_in = testData4[204];
@(posedge clk);
#1;data_in = testData4[205];
@(posedge clk);
#1;data_in = testData4[206];
@(posedge clk);
#1;data_in = testData4[207];
@(posedge clk);
#1;data_in = testData4[208];
@(posedge clk);
#1;data_in = testData4[209];
@(posedge clk);
#1;data_in = testData4[210];
@(posedge clk);
#1;data_in = testData4[211];
@(posedge clk);
#1;data_in = testData4[212];
@(posedge clk);
#1;data_in = testData4[213];
@(posedge clk);
#1;data_in = testData4[214];
@(posedge clk);
#1;data_in = testData4[215];
@(posedge clk);
#1;data_in = testData4[216];
@(posedge clk);
#1;data_in = testData4[217];
@(posedge clk);
#1;data_in = testData4[218];
@(posedge clk);
#1;data_in = testData4[219];
@(posedge clk);
#1;data_in = testData4[220];
@(posedge clk);
#1;data_in = testData4[221];
@(posedge clk);
#1;data_in = testData4[222];
@(posedge clk);
#1;data_in = testData4[223];
@(posedge clk);
#1;data_in = testData4[224];
@(posedge clk);
#1;data_in = testData4[225];
@(posedge clk);
#1;data_in = testData4[226];
@(posedge clk);
#1;data_in = testData4[227];
@(posedge clk);
#1;data_in = testData4[228];
@(posedge clk);
#1;data_in = testData4[229];
@(posedge clk);
#1;data_in = testData4[230];
@(posedge clk);
#1;data_in = testData4[231];
@(posedge clk);
#1;data_in = testData4[232];
@(posedge clk);
#1;data_in = testData4[233];
@(posedge clk);
#1;data_in = testData4[234];
@(posedge clk);
#1;data_in = testData4[235];
@(posedge clk);
#1;data_in = testData4[236];
@(posedge clk);
#1;data_in = testData4[237];
@(posedge clk);
#1;data_in = testData4[238];
@(posedge clk);
#1;data_in = testData4[239];
@(posedge clk);
#1;data_in = testData4[240];
@(posedge clk);
#1;data_in = testData4[241];
@(posedge clk);
#1;data_in = testData4[242];
@(posedge clk);
#1;data_in = testData4[243];
@(posedge clk);
#1;data_in = testData4[244];
@(posedge clk);
#1;data_in = testData4[245];
@(posedge clk);
#1;data_in = testData4[246];
@(posedge clk);
#1;data_in = testData4[247];
@(posedge clk);
#1;data_in = testData4[248];
@(posedge clk);
#1;data_in = testData4[249];
@(posedge clk);
#1;data_in = testData4[250];
@(posedge clk);
#1;data_in = testData4[251];
@(posedge clk);
#1;data_in = testData4[252];
@(posedge clk);
#1;data_in = testData4[253];
@(posedge clk);
#1;data_in = testData4[254];
@(posedge clk);
#1;data_in = testData4[255];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData4[256]; 
@(posedge clk);
#1;data_in = testData4[257];
@(posedge clk);
#1;data_in = testData4[258];
@(posedge clk);
#1;data_in = testData4[259];
@(posedge clk);
#1;data_in = testData4[260];
@(posedge clk);
#1;data_in = testData4[261];
@(posedge clk);
#1;data_in = testData4[262];
@(posedge clk);
#1;data_in = testData4[263];
@(posedge clk);
#1;data_in = testData4[264];
@(posedge clk);
#1;data_in = testData4[265];
@(posedge clk);
#1;data_in = testData4[266];
@(posedge clk);
#1;data_in = testData4[267];
@(posedge clk);
#1;data_in = testData4[268];
@(posedge clk);
#1;data_in = testData4[269];
@(posedge clk);
#1;data_in = testData4[270];
@(posedge clk);
#1;data_in = testData4[271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[272]; 
@(posedge clk);
#1;data_in = testData4[273];
@(posedge clk);
#1;data_in = testData4[274];
@(posedge clk);
#1;data_in = testData4[275];
@(posedge clk);
#1;data_in = testData4[276];
@(posedge clk);
#1;data_in = testData4[277];
@(posedge clk);
#1;data_in = testData4[278];
@(posedge clk);
#1;data_in = testData4[279];
@(posedge clk);
#1;data_in = testData4[280];
@(posedge clk);
#1;data_in = testData4[281];
@(posedge clk);
#1;data_in = testData4[282];
@(posedge clk);
#1;data_in = testData4[283];
@(posedge clk);
#1;data_in = testData4[284];
@(posedge clk);
#1;data_in = testData4[285];
@(posedge clk);
#1;data_in = testData4[286];
@(posedge clk);
#1;data_in = testData4[287];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[288]; 
@(posedge clk);
#1;data_in = testData4[289];
@(posedge clk);
#1;data_in = testData4[290];
@(posedge clk);
#1;data_in = testData4[291];
@(posedge clk);
#1;data_in = testData4[292];
@(posedge clk);
#1;data_in = testData4[293];
@(posedge clk);
#1;data_in = testData4[294];
@(posedge clk);
#1;data_in = testData4[295];
@(posedge clk);
#1;data_in = testData4[296];
@(posedge clk);
#1;data_in = testData4[297];
@(posedge clk);
#1;data_in = testData4[298];
@(posedge clk);
#1;data_in = testData4[299];
@(posedge clk);
#1;data_in = testData4[300];
@(posedge clk);
#1;data_in = testData4[301];
@(posedge clk);
#1;data_in = testData4[302];
@(posedge clk);
#1;data_in = testData4[303];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[304]; 
@(posedge clk);
#1;data_in = testData4[305];
@(posedge clk);
#1;data_in = testData4[306];
@(posedge clk);
#1;data_in = testData4[307];
@(posedge clk);
#1;data_in = testData4[308];
@(posedge clk);
#1;data_in = testData4[309];
@(posedge clk);
#1;data_in = testData4[310];
@(posedge clk);
#1;data_in = testData4[311];
@(posedge clk);
#1;data_in = testData4[312];
@(posedge clk);
#1;data_in = testData4[313];
@(posedge clk);
#1;data_in = testData4[314];
@(posedge clk);
#1;data_in = testData4[315];
@(posedge clk);
#1;data_in = testData4[316];
@(posedge clk);
#1;data_in = testData4[317];
@(posedge clk);
#1;data_in = testData4[318];
@(posedge clk);
#1;data_in = testData4[319];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[320]; 
@(posedge clk);
#1;data_in = testData4[321];
@(posedge clk);
#1;data_in = testData4[322];
@(posedge clk);
#1;data_in = testData4[323];
@(posedge clk);
#1;data_in = testData4[324];
@(posedge clk);
#1;data_in = testData4[325];
@(posedge clk);
#1;data_in = testData4[326];
@(posedge clk);
#1;data_in = testData4[327];
@(posedge clk);
#1;data_in = testData4[328];
@(posedge clk);
#1;data_in = testData4[329];
@(posedge clk);
#1;data_in = testData4[330];
@(posedge clk);
#1;data_in = testData4[331];
@(posedge clk);
#1;data_in = testData4[332];
@(posedge clk);
#1;data_in = testData4[333];
@(posedge clk);
#1;data_in = testData4[334];
@(posedge clk);
#1;data_in = testData4[335];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[336]; 
@(posedge clk);
#1;data_in = testData4[337];
@(posedge clk);
#1;data_in = testData4[338];
@(posedge clk);
#1;data_in = testData4[339];
@(posedge clk);
#1;data_in = testData4[340];
@(posedge clk);
#1;data_in = testData4[341];
@(posedge clk);
#1;data_in = testData4[342];
@(posedge clk);
#1;data_in = testData4[343];
@(posedge clk);
#1;data_in = testData4[344];
@(posedge clk);
#1;data_in = testData4[345];
@(posedge clk);
#1;data_in = testData4[346];
@(posedge clk);
#1;data_in = testData4[347];
@(posedge clk);
#1;data_in = testData4[348];
@(posedge clk);
#1;data_in = testData4[349];
@(posedge clk);
#1;data_in = testData4[350];
@(posedge clk);
#1;data_in = testData4[351];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[352]; 
@(posedge clk);
#1;data_in = testData4[353];
@(posedge clk);
#1;data_in = testData4[354];
@(posedge clk);
#1;data_in = testData4[355];
@(posedge clk);
#1;data_in = testData4[356];
@(posedge clk);
#1;data_in = testData4[357];
@(posedge clk);
#1;data_in = testData4[358];
@(posedge clk);
#1;data_in = testData4[359];
@(posedge clk);
#1;data_in = testData4[360];
@(posedge clk);
#1;data_in = testData4[361];
@(posedge clk);
#1;data_in = testData4[362];
@(posedge clk);
#1;data_in = testData4[363];
@(posedge clk);
#1;data_in = testData4[364];
@(posedge clk);
#1;data_in = testData4[365];
@(posedge clk);
#1;data_in = testData4[366];
@(posedge clk);
#1;data_in = testData4[367];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[368]; 
@(posedge clk);
#1;data_in = testData4[369];
@(posedge clk);
#1;data_in = testData4[370];
@(posedge clk);
#1;data_in = testData4[371];
@(posedge clk);
#1;data_in = testData4[372];
@(posedge clk);
#1;data_in = testData4[373];
@(posedge clk);
#1;data_in = testData4[374];
@(posedge clk);
#1;data_in = testData4[375];
@(posedge clk);
#1;data_in = testData4[376];
@(posedge clk);
#1;data_in = testData4[377];
@(posedge clk);
#1;data_in = testData4[378];
@(posedge clk);
#1;data_in = testData4[379];
@(posedge clk);
#1;data_in = testData4[380];
@(posedge clk);
#1;data_in = testData4[381];
@(posedge clk);
#1;data_in = testData4[382];
@(posedge clk);
#1;data_in = testData4[383];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[384]; 
@(posedge clk);
#1;data_in = testData4[385];
@(posedge clk);
#1;data_in = testData4[386];
@(posedge clk);
#1;data_in = testData4[387];
@(posedge clk);
#1;data_in = testData4[388];
@(posedge clk);
#1;data_in = testData4[389];
@(posedge clk);
#1;data_in = testData4[390];
@(posedge clk);
#1;data_in = testData4[391];
@(posedge clk);
#1;data_in = testData4[392];
@(posedge clk);
#1;data_in = testData4[393];
@(posedge clk);
#1;data_in = testData4[394];
@(posedge clk);
#1;data_in = testData4[395];
@(posedge clk);
#1;data_in = testData4[396];
@(posedge clk);
#1;data_in = testData4[397];
@(posedge clk);
#1;data_in = testData4[398];
@(posedge clk);
#1;data_in = testData4[399];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[400]; 
@(posedge clk);
#1;data_in = testData4[401];
@(posedge clk);
#1;data_in = testData4[402];
@(posedge clk);
#1;data_in = testData4[403];
@(posedge clk);
#1;data_in = testData4[404];
@(posedge clk);
#1;data_in = testData4[405];
@(posedge clk);
#1;data_in = testData4[406];
@(posedge clk);
#1;data_in = testData4[407];
@(posedge clk);
#1;data_in = testData4[408];
@(posedge clk);
#1;data_in = testData4[409];
@(posedge clk);
#1;data_in = testData4[410];
@(posedge clk);
#1;data_in = testData4[411];
@(posedge clk);
#1;data_in = testData4[412];
@(posedge clk);
#1;data_in = testData4[413];
@(posedge clk);
#1;data_in = testData4[414];
@(posedge clk);
#1;data_in = testData4[415];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[416]; 
@(posedge clk);
#1;data_in = testData4[417];
@(posedge clk);
#1;data_in = testData4[418];
@(posedge clk);
#1;data_in = testData4[419];
@(posedge clk);
#1;data_in = testData4[420];
@(posedge clk);
#1;data_in = testData4[421];
@(posedge clk);
#1;data_in = testData4[422];
@(posedge clk);
#1;data_in = testData4[423];
@(posedge clk);
#1;data_in = testData4[424];
@(posedge clk);
#1;data_in = testData4[425];
@(posedge clk);
#1;data_in = testData4[426];
@(posedge clk);
#1;data_in = testData4[427];
@(posedge clk);
#1;data_in = testData4[428];
@(posedge clk);
#1;data_in = testData4[429];
@(posedge clk);
#1;data_in = testData4[430];
@(posedge clk);
#1;data_in = testData4[431];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[432]; 
@(posedge clk);
#1;data_in = testData4[433];
@(posedge clk);
#1;data_in = testData4[434];
@(posedge clk);
#1;data_in = testData4[435];
@(posedge clk);
#1;data_in = testData4[436];
@(posedge clk);
#1;data_in = testData4[437];
@(posedge clk);
#1;data_in = testData4[438];
@(posedge clk);
#1;data_in = testData4[439];
@(posedge clk);
#1;data_in = testData4[440];
@(posedge clk);
#1;data_in = testData4[441];
@(posedge clk);
#1;data_in = testData4[442];
@(posedge clk);
#1;data_in = testData4[443];
@(posedge clk);
#1;data_in = testData4[444];
@(posedge clk);
#1;data_in = testData4[445];
@(posedge clk);
#1;data_in = testData4[446];
@(posedge clk);
#1;data_in = testData4[447];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[448]; 
@(posedge clk);
#1;data_in = testData4[449];
@(posedge clk);
#1;data_in = testData4[450];
@(posedge clk);
#1;data_in = testData4[451];
@(posedge clk);
#1;data_in = testData4[452];
@(posedge clk);
#1;data_in = testData4[453];
@(posedge clk);
#1;data_in = testData4[454];
@(posedge clk);
#1;data_in = testData4[455];
@(posedge clk);
#1;data_in = testData4[456];
@(posedge clk);
#1;data_in = testData4[457];
@(posedge clk);
#1;data_in = testData4[458];
@(posedge clk);
#1;data_in = testData4[459];
@(posedge clk);
#1;data_in = testData4[460];
@(posedge clk);
#1;data_in = testData4[461];
@(posedge clk);
#1;data_in = testData4[462];
@(posedge clk);
#1;data_in = testData4[463];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[464]; 
@(posedge clk);
#1;data_in = testData4[465];
@(posedge clk);
#1;data_in = testData4[466];
@(posedge clk);
#1;data_in = testData4[467];
@(posedge clk);
#1;data_in = testData4[468];
@(posedge clk);
#1;data_in = testData4[469];
@(posedge clk);
#1;data_in = testData4[470];
@(posedge clk);
#1;data_in = testData4[471];
@(posedge clk);
#1;data_in = testData4[472];
@(posedge clk);
#1;data_in = testData4[473];
@(posedge clk);
#1;data_in = testData4[474];
@(posedge clk);
#1;data_in = testData4[475];
@(posedge clk);
#1;data_in = testData4[476];
@(posedge clk);
#1;data_in = testData4[477];
@(posedge clk);
#1;data_in = testData4[478];
@(posedge clk);
#1;data_in = testData4[479];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[480]; 
@(posedge clk);
#1;data_in = testData4[481];
@(posedge clk);
#1;data_in = testData4[482];
@(posedge clk);
#1;data_in = testData4[483];
@(posedge clk);
#1;data_in = testData4[484];
@(posedge clk);
#1;data_in = testData4[485];
@(posedge clk);
#1;data_in = testData4[486];
@(posedge clk);
#1;data_in = testData4[487];
@(posedge clk);
#1;data_in = testData4[488];
@(posedge clk);
#1;data_in = testData4[489];
@(posedge clk);
#1;data_in = testData4[490];
@(posedge clk);
#1;data_in = testData4[491];
@(posedge clk);
#1;data_in = testData4[492];
@(posedge clk);
#1;data_in = testData4[493];
@(posedge clk);
#1;data_in = testData4[494];
@(posedge clk);
#1;data_in = testData4[495];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[496]; 
@(posedge clk);
#1;data_in = testData4[497];
@(posedge clk);
#1;data_in = testData4[498];
@(posedge clk);
#1;data_in = testData4[499];
@(posedge clk);
#1;data_in = testData4[500];
@(posedge clk);
#1;data_in = testData4[501];
@(posedge clk);
#1;data_in = testData4[502];
@(posedge clk);
#1;data_in = testData4[503];
@(posedge clk);
#1;data_in = testData4[504];
@(posedge clk);
#1;data_in = testData4[505];
@(posedge clk);
#1;data_in = testData4[506];
@(posedge clk);
#1;data_in = testData4[507];
@(posedge clk);
#1;data_in = testData4[508];
@(posedge clk);
#1;data_in = testData4[509];
@(posedge clk);
#1;data_in = testData4[510];
@(posedge clk);
#1;data_in = testData4[511];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[512]; 
@(posedge clk);
#1;data_in = testData4[513];
@(posedge clk);
#1;data_in = testData4[514];
@(posedge clk);
#1;data_in = testData4[515];
@(posedge clk);
#1;data_in = testData4[516];
@(posedge clk);
#1;data_in = testData4[517];
@(posedge clk);
#1;data_in = testData4[518];
@(posedge clk);
#1;data_in = testData4[519];
@(posedge clk);
#1;data_in = testData4[520];
@(posedge clk);
#1;data_in = testData4[521];
@(posedge clk);
#1;data_in = testData4[522];
@(posedge clk);
#1;data_in = testData4[523];
@(posedge clk);
#1;data_in = testData4[524];
@(posedge clk);
#1;data_in = testData4[525];
@(posedge clk);
#1;data_in = testData4[526];
@(posedge clk);
#1;data_in = testData4[527];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[528]; 
@(posedge clk);
#1;data_in = testData4[529];
@(posedge clk);
#1;data_in = testData4[530];
@(posedge clk);
#1;data_in = testData4[531];
@(posedge clk);
#1;data_in = testData4[532];
@(posedge clk);
#1;data_in = testData4[533];
@(posedge clk);
#1;data_in = testData4[534];
@(posedge clk);
#1;data_in = testData4[535];
@(posedge clk);
#1;data_in = testData4[536];
@(posedge clk);
#1;data_in = testData4[537];
@(posedge clk);
#1;data_in = testData4[538];
@(posedge clk);
#1;data_in = testData4[539];
@(posedge clk);
#1;data_in = testData4[540];
@(posedge clk);
#1;data_in = testData4[541];
@(posedge clk);
#1;data_in = testData4[542];
@(posedge clk);
#1;data_in = testData4[543];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[544]; 
@(posedge clk);
#1;data_in = testData4[545];
@(posedge clk);
#1;data_in = testData4[546];
@(posedge clk);
#1;data_in = testData4[547];
@(posedge clk);
#1;data_in = testData4[548];
@(posedge clk);
#1;data_in = testData4[549];
@(posedge clk);
#1;data_in = testData4[550];
@(posedge clk);
#1;data_in = testData4[551];
@(posedge clk);
#1;data_in = testData4[552];
@(posedge clk);
#1;data_in = testData4[553];
@(posedge clk);
#1;data_in = testData4[554];
@(posedge clk);
#1;data_in = testData4[555];
@(posedge clk);
#1;data_in = testData4[556];
@(posedge clk);
#1;data_in = testData4[557];
@(posedge clk);
#1;data_in = testData4[558];
@(posedge clk);
#1;data_in = testData4[559];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[560]; 
@(posedge clk);
#1;data_in = testData4[561];
@(posedge clk);
#1;data_in = testData4[562];
@(posedge clk);
#1;data_in = testData4[563];
@(posedge clk);
#1;data_in = testData4[564];
@(posedge clk);
#1;data_in = testData4[565];
@(posedge clk);
#1;data_in = testData4[566];
@(posedge clk);
#1;data_in = testData4[567];
@(posedge clk);
#1;data_in = testData4[568];
@(posedge clk);
#1;data_in = testData4[569];
@(posedge clk);
#1;data_in = testData4[570];
@(posedge clk);
#1;data_in = testData4[571];
@(posedge clk);
#1;data_in = testData4[572];
@(posedge clk);
#1;data_in = testData4[573];
@(posedge clk);
#1;data_in = testData4[574];
@(posedge clk);
#1;data_in = testData4[575];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[576]; 
@(posedge clk);
#1;data_in = testData4[577];
@(posedge clk);
#1;data_in = testData4[578];
@(posedge clk);
#1;data_in = testData4[579];
@(posedge clk);
#1;data_in = testData4[580];
@(posedge clk);
#1;data_in = testData4[581];
@(posedge clk);
#1;data_in = testData4[582];
@(posedge clk);
#1;data_in = testData4[583];
@(posedge clk);
#1;data_in = testData4[584];
@(posedge clk);
#1;data_in = testData4[585];
@(posedge clk);
#1;data_in = testData4[586];
@(posedge clk);
#1;data_in = testData4[587];
@(posedge clk);
#1;data_in = testData4[588];
@(posedge clk);
#1;data_in = testData4[589];
@(posedge clk);
#1;data_in = testData4[590];
@(posedge clk);
#1;data_in = testData4[591];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[592]; 
@(posedge clk);
#1;data_in = testData4[593];
@(posedge clk);
#1;data_in = testData4[594];
@(posedge clk);
#1;data_in = testData4[595];
@(posedge clk);
#1;data_in = testData4[596];
@(posedge clk);
#1;data_in = testData4[597];
@(posedge clk);
#1;data_in = testData4[598];
@(posedge clk);
#1;data_in = testData4[599];
@(posedge clk);
#1;data_in = testData4[600];
@(posedge clk);
#1;data_in = testData4[601];
@(posedge clk);
#1;data_in = testData4[602];
@(posedge clk);
#1;data_in = testData4[603];
@(posedge clk);
#1;data_in = testData4[604];
@(posedge clk);
#1;data_in = testData4[605];
@(posedge clk);
#1;data_in = testData4[606];
@(posedge clk);
#1;data_in = testData4[607];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[608]; 
@(posedge clk);
#1;data_in = testData4[609];
@(posedge clk);
#1;data_in = testData4[610];
@(posedge clk);
#1;data_in = testData4[611];
@(posedge clk);
#1;data_in = testData4[612];
@(posedge clk);
#1;data_in = testData4[613];
@(posedge clk);
#1;data_in = testData4[614];
@(posedge clk);
#1;data_in = testData4[615];
@(posedge clk);
#1;data_in = testData4[616];
@(posedge clk);
#1;data_in = testData4[617];
@(posedge clk);
#1;data_in = testData4[618];
@(posedge clk);
#1;data_in = testData4[619];
@(posedge clk);
#1;data_in = testData4[620];
@(posedge clk);
#1;data_in = testData4[621];
@(posedge clk);
#1;data_in = testData4[622];
@(posedge clk);
#1;data_in = testData4[623];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[624]; 
@(posedge clk);
#1;data_in = testData4[625];
@(posedge clk);
#1;data_in = testData4[626];
@(posedge clk);
#1;data_in = testData4[627];
@(posedge clk);
#1;data_in = testData4[628];
@(posedge clk);
#1;data_in = testData4[629];
@(posedge clk);
#1;data_in = testData4[630];
@(posedge clk);
#1;data_in = testData4[631];
@(posedge clk);
#1;data_in = testData4[632];
@(posedge clk);
#1;data_in = testData4[633];
@(posedge clk);
#1;data_in = testData4[634];
@(posedge clk);
#1;data_in = testData4[635];
@(posedge clk);
#1;data_in = testData4[636];
@(posedge clk);
#1;data_in = testData4[637];
@(posedge clk);
#1;data_in = testData4[638];
@(posedge clk);
#1;data_in = testData4[639];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[640]; 
@(posedge clk);
#1;data_in = testData4[641];
@(posedge clk);
#1;data_in = testData4[642];
@(posedge clk);
#1;data_in = testData4[643];
@(posedge clk);
#1;data_in = testData4[644];
@(posedge clk);
#1;data_in = testData4[645];
@(posedge clk);
#1;data_in = testData4[646];
@(posedge clk);
#1;data_in = testData4[647];
@(posedge clk);
#1;data_in = testData4[648];
@(posedge clk);
#1;data_in = testData4[649];
@(posedge clk);
#1;data_in = testData4[650];
@(posedge clk);
#1;data_in = testData4[651];
@(posedge clk);
#1;data_in = testData4[652];
@(posedge clk);
#1;data_in = testData4[653];
@(posedge clk);
#1;data_in = testData4[654];
@(posedge clk);
#1;data_in = testData4[655];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[656]; 
@(posedge clk);
#1;data_in = testData4[657];
@(posedge clk);
#1;data_in = testData4[658];
@(posedge clk);
#1;data_in = testData4[659];
@(posedge clk);
#1;data_in = testData4[660];
@(posedge clk);
#1;data_in = testData4[661];
@(posedge clk);
#1;data_in = testData4[662];
@(posedge clk);
#1;data_in = testData4[663];
@(posedge clk);
#1;data_in = testData4[664];
@(posedge clk);
#1;data_in = testData4[665];
@(posedge clk);
#1;data_in = testData4[666];
@(posedge clk);
#1;data_in = testData4[667];
@(posedge clk);
#1;data_in = testData4[668];
@(posedge clk);
#1;data_in = testData4[669];
@(posedge clk);
#1;data_in = testData4[670];
@(posedge clk);
#1;data_in = testData4[671];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[672]; 
@(posedge clk);
#1;data_in = testData4[673];
@(posedge clk);
#1;data_in = testData4[674];
@(posedge clk);
#1;data_in = testData4[675];
@(posedge clk);
#1;data_in = testData4[676];
@(posedge clk);
#1;data_in = testData4[677];
@(posedge clk);
#1;data_in = testData4[678];
@(posedge clk);
#1;data_in = testData4[679];
@(posedge clk);
#1;data_in = testData4[680];
@(posedge clk);
#1;data_in = testData4[681];
@(posedge clk);
#1;data_in = testData4[682];
@(posedge clk);
#1;data_in = testData4[683];
@(posedge clk);
#1;data_in = testData4[684];
@(posedge clk);
#1;data_in = testData4[685];
@(posedge clk);
#1;data_in = testData4[686];
@(posedge clk);
#1;data_in = testData4[687];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[688]; 
@(posedge clk);
#1;data_in = testData4[689];
@(posedge clk);
#1;data_in = testData4[690];
@(posedge clk);
#1;data_in = testData4[691];
@(posedge clk);
#1;data_in = testData4[692];
@(posedge clk);
#1;data_in = testData4[693];
@(posedge clk);
#1;data_in = testData4[694];
@(posedge clk);
#1;data_in = testData4[695];
@(posedge clk);
#1;data_in = testData4[696];
@(posedge clk);
#1;data_in = testData4[697];
@(posedge clk);
#1;data_in = testData4[698];
@(posedge clk);
#1;data_in = testData4[699];
@(posedge clk);
#1;data_in = testData4[700];
@(posedge clk);
#1;data_in = testData4[701];
@(posedge clk);
#1;data_in = testData4[702];
@(posedge clk);
#1;data_in = testData4[703];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[704]; 
@(posedge clk);
#1;data_in = testData4[705];
@(posedge clk);
#1;data_in = testData4[706];
@(posedge clk);
#1;data_in = testData4[707];
@(posedge clk);
#1;data_in = testData4[708];
@(posedge clk);
#1;data_in = testData4[709];
@(posedge clk);
#1;data_in = testData4[710];
@(posedge clk);
#1;data_in = testData4[711];
@(posedge clk);
#1;data_in = testData4[712];
@(posedge clk);
#1;data_in = testData4[713];
@(posedge clk);
#1;data_in = testData4[714];
@(posedge clk);
#1;data_in = testData4[715];
@(posedge clk);
#1;data_in = testData4[716];
@(posedge clk);
#1;data_in = testData4[717];
@(posedge clk);
#1;data_in = testData4[718];
@(posedge clk);
#1;data_in = testData4[719];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[720]; 
@(posedge clk);
#1;data_in = testData4[721];
@(posedge clk);
#1;data_in = testData4[722];
@(posedge clk);
#1;data_in = testData4[723];
@(posedge clk);
#1;data_in = testData4[724];
@(posedge clk);
#1;data_in = testData4[725];
@(posedge clk);
#1;data_in = testData4[726];
@(posedge clk);
#1;data_in = testData4[727];
@(posedge clk);
#1;data_in = testData4[728];
@(posedge clk);
#1;data_in = testData4[729];
@(posedge clk);
#1;data_in = testData4[730];
@(posedge clk);
#1;data_in = testData4[731];
@(posedge clk);
#1;data_in = testData4[732];
@(posedge clk);
#1;data_in = testData4[733];
@(posedge clk);
#1;data_in = testData4[734];
@(posedge clk);
#1;data_in = testData4[735];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[736]; 
@(posedge clk);
#1;data_in = testData4[737];
@(posedge clk);
#1;data_in = testData4[738];
@(posedge clk);
#1;data_in = testData4[739];
@(posedge clk);
#1;data_in = testData4[740];
@(posedge clk);
#1;data_in = testData4[741];
@(posedge clk);
#1;data_in = testData4[742];
@(posedge clk);
#1;data_in = testData4[743];
@(posedge clk);
#1;data_in = testData4[744];
@(posedge clk);
#1;data_in = testData4[745];
@(posedge clk);
#1;data_in = testData4[746];
@(posedge clk);
#1;data_in = testData4[747];
@(posedge clk);
#1;data_in = testData4[748];
@(posedge clk);
#1;data_in = testData4[749];
@(posedge clk);
#1;data_in = testData4[750];
@(posedge clk);
#1;data_in = testData4[751];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[752]; 
@(posedge clk);
#1;data_in = testData4[753];
@(posedge clk);
#1;data_in = testData4[754];
@(posedge clk);
#1;data_in = testData4[755];
@(posedge clk);
#1;data_in = testData4[756];
@(posedge clk);
#1;data_in = testData4[757];
@(posedge clk);
#1;data_in = testData4[758];
@(posedge clk);
#1;data_in = testData4[759];
@(posedge clk);
#1;data_in = testData4[760];
@(posedge clk);
#1;data_in = testData4[761];
@(posedge clk);
#1;data_in = testData4[762];
@(posedge clk);
#1;data_in = testData4[763];
@(posedge clk);
#1;data_in = testData4[764];
@(posedge clk);
#1;data_in = testData4[765];
@(posedge clk);
#1;data_in = testData4[766];
@(posedge clk);
#1;data_in = testData4[767];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[768]; 
@(posedge clk);
#1;data_in = testData4[769];
@(posedge clk);
#1;data_in = testData4[770];
@(posedge clk);
#1;data_in = testData4[771];
@(posedge clk);
#1;data_in = testData4[772];
@(posedge clk);
#1;data_in = testData4[773];
@(posedge clk);
#1;data_in = testData4[774];
@(posedge clk);
#1;data_in = testData4[775];
@(posedge clk);
#1;data_in = testData4[776];
@(posedge clk);
#1;data_in = testData4[777];
@(posedge clk);
#1;data_in = testData4[778];
@(posedge clk);
#1;data_in = testData4[779];
@(posedge clk);
#1;data_in = testData4[780];
@(posedge clk);
#1;data_in = testData4[781];
@(posedge clk);
#1;data_in = testData4[782];
@(posedge clk);
#1;data_in = testData4[783];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[784]; 
@(posedge clk);
#1;data_in = testData4[785];
@(posedge clk);
#1;data_in = testData4[786];
@(posedge clk);
#1;data_in = testData4[787];
@(posedge clk);
#1;data_in = testData4[788];
@(posedge clk);
#1;data_in = testData4[789];
@(posedge clk);
#1;data_in = testData4[790];
@(posedge clk);
#1;data_in = testData4[791];
@(posedge clk);
#1;data_in = testData4[792];
@(posedge clk);
#1;data_in = testData4[793];
@(posedge clk);
#1;data_in = testData4[794];
@(posedge clk);
#1;data_in = testData4[795];
@(posedge clk);
#1;data_in = testData4[796];
@(posedge clk);
#1;data_in = testData4[797];
@(posedge clk);
#1;data_in = testData4[798];
@(posedge clk);
#1;data_in = testData4[799];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[800]; 
@(posedge clk);
#1;data_in = testData4[801];
@(posedge clk);
#1;data_in = testData4[802];
@(posedge clk);
#1;data_in = testData4[803];
@(posedge clk);
#1;data_in = testData4[804];
@(posedge clk);
#1;data_in = testData4[805];
@(posedge clk);
#1;data_in = testData4[806];
@(posedge clk);
#1;data_in = testData4[807];
@(posedge clk);
#1;data_in = testData4[808];
@(posedge clk);
#1;data_in = testData4[809];
@(posedge clk);
#1;data_in = testData4[810];
@(posedge clk);
#1;data_in = testData4[811];
@(posedge clk);
#1;data_in = testData4[812];
@(posedge clk);
#1;data_in = testData4[813];
@(posedge clk);
#1;data_in = testData4[814];
@(posedge clk);
#1;data_in = testData4[815];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[816]; 
@(posedge clk);
#1;data_in = testData4[817];
@(posedge clk);
#1;data_in = testData4[818];
@(posedge clk);
#1;data_in = testData4[819];
@(posedge clk);
#1;data_in = testData4[820];
@(posedge clk);
#1;data_in = testData4[821];
@(posedge clk);
#1;data_in = testData4[822];
@(posedge clk);
#1;data_in = testData4[823];
@(posedge clk);
#1;data_in = testData4[824];
@(posedge clk);
#1;data_in = testData4[825];
@(posedge clk);
#1;data_in = testData4[826];
@(posedge clk);
#1;data_in = testData4[827];
@(posedge clk);
#1;data_in = testData4[828];
@(posedge clk);
#1;data_in = testData4[829];
@(posedge clk);
#1;data_in = testData4[830];
@(posedge clk);
#1;data_in = testData4[831];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[832]; 
@(posedge clk);
#1;data_in = testData4[833];
@(posedge clk);
#1;data_in = testData4[834];
@(posedge clk);
#1;data_in = testData4[835];
@(posedge clk);
#1;data_in = testData4[836];
@(posedge clk);
#1;data_in = testData4[837];
@(posedge clk);
#1;data_in = testData4[838];
@(posedge clk);
#1;data_in = testData4[839];
@(posedge clk);
#1;data_in = testData4[840];
@(posedge clk);
#1;data_in = testData4[841];
@(posedge clk);
#1;data_in = testData4[842];
@(posedge clk);
#1;data_in = testData4[843];
@(posedge clk);
#1;data_in = testData4[844];
@(posedge clk);
#1;data_in = testData4[845];
@(posedge clk);
#1;data_in = testData4[846];
@(posedge clk);
#1;data_in = testData4[847];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[848]; 
@(posedge clk);
#1;data_in = testData4[849];
@(posedge clk);
#1;data_in = testData4[850];
@(posedge clk);
#1;data_in = testData4[851];
@(posedge clk);
#1;data_in = testData4[852];
@(posedge clk);
#1;data_in = testData4[853];
@(posedge clk);
#1;data_in = testData4[854];
@(posedge clk);
#1;data_in = testData4[855];
@(posedge clk);
#1;data_in = testData4[856];
@(posedge clk);
#1;data_in = testData4[857];
@(posedge clk);
#1;data_in = testData4[858];
@(posedge clk);
#1;data_in = testData4[859];
@(posedge clk);
#1;data_in = testData4[860];
@(posedge clk);
#1;data_in = testData4[861];
@(posedge clk);
#1;data_in = testData4[862];
@(posedge clk);
#1;data_in = testData4[863];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[864]; 
@(posedge clk);
#1;data_in = testData4[865];
@(posedge clk);
#1;data_in = testData4[866];
@(posedge clk);
#1;data_in = testData4[867];
@(posedge clk);
#1;data_in = testData4[868];
@(posedge clk);
#1;data_in = testData4[869];
@(posedge clk);
#1;data_in = testData4[870];
@(posedge clk);
#1;data_in = testData4[871];
@(posedge clk);
#1;data_in = testData4[872];
@(posedge clk);
#1;data_in = testData4[873];
@(posedge clk);
#1;data_in = testData4[874];
@(posedge clk);
#1;data_in = testData4[875];
@(posedge clk);
#1;data_in = testData4[876];
@(posedge clk);
#1;data_in = testData4[877];
@(posedge clk);
#1;data_in = testData4[878];
@(posedge clk);
#1;data_in = testData4[879];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[880]; 
@(posedge clk);
#1;data_in = testData4[881];
@(posedge clk);
#1;data_in = testData4[882];
@(posedge clk);
#1;data_in = testData4[883];
@(posedge clk);
#1;data_in = testData4[884];
@(posedge clk);
#1;data_in = testData4[885];
@(posedge clk);
#1;data_in = testData4[886];
@(posedge clk);
#1;data_in = testData4[887];
@(posedge clk);
#1;data_in = testData4[888];
@(posedge clk);
#1;data_in = testData4[889];
@(posedge clk);
#1;data_in = testData4[890];
@(posedge clk);
#1;data_in = testData4[891];
@(posedge clk);
#1;data_in = testData4[892];
@(posedge clk);
#1;data_in = testData4[893];
@(posedge clk);
#1;data_in = testData4[894];
@(posedge clk);
#1;data_in = testData4[895];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[896]; 
@(posedge clk);
#1;data_in = testData4[897];
@(posedge clk);
#1;data_in = testData4[898];
@(posedge clk);
#1;data_in = testData4[899];
@(posedge clk);
#1;data_in = testData4[900];
@(posedge clk);
#1;data_in = testData4[901];
@(posedge clk);
#1;data_in = testData4[902];
@(posedge clk);
#1;data_in = testData4[903];
@(posedge clk);
#1;data_in = testData4[904];
@(posedge clk);
#1;data_in = testData4[905];
@(posedge clk);
#1;data_in = testData4[906];
@(posedge clk);
#1;data_in = testData4[907];
@(posedge clk);
#1;data_in = testData4[908];
@(posedge clk);
#1;data_in = testData4[909];
@(posedge clk);
#1;data_in = testData4[910];
@(posedge clk);
#1;data_in = testData4[911];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[912]; 
@(posedge clk);
#1;data_in = testData4[913];
@(posedge clk);
#1;data_in = testData4[914];
@(posedge clk);
#1;data_in = testData4[915];
@(posedge clk);
#1;data_in = testData4[916];
@(posedge clk);
#1;data_in = testData4[917];
@(posedge clk);
#1;data_in = testData4[918];
@(posedge clk);
#1;data_in = testData4[919];
@(posedge clk);
#1;data_in = testData4[920];
@(posedge clk);
#1;data_in = testData4[921];
@(posedge clk);
#1;data_in = testData4[922];
@(posedge clk);
#1;data_in = testData4[923];
@(posedge clk);
#1;data_in = testData4[924];
@(posedge clk);
#1;data_in = testData4[925];
@(posedge clk);
#1;data_in = testData4[926];
@(posedge clk);
#1;data_in = testData4[927];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[928]; 
@(posedge clk);
#1;data_in = testData4[929];
@(posedge clk);
#1;data_in = testData4[930];
@(posedge clk);
#1;data_in = testData4[931];
@(posedge clk);
#1;data_in = testData4[932];
@(posedge clk);
#1;data_in = testData4[933];
@(posedge clk);
#1;data_in = testData4[934];
@(posedge clk);
#1;data_in = testData4[935];
@(posedge clk);
#1;data_in = testData4[936];
@(posedge clk);
#1;data_in = testData4[937];
@(posedge clk);
#1;data_in = testData4[938];
@(posedge clk);
#1;data_in = testData4[939];
@(posedge clk);
#1;data_in = testData4[940];
@(posedge clk);
#1;data_in = testData4[941];
@(posedge clk);
#1;data_in = testData4[942];
@(posedge clk);
#1;data_in = testData4[943];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[944]; 
@(posedge clk);
#1;data_in = testData4[945];
@(posedge clk);
#1;data_in = testData4[946];
@(posedge clk);
#1;data_in = testData4[947];
@(posedge clk);
#1;data_in = testData4[948];
@(posedge clk);
#1;data_in = testData4[949];
@(posedge clk);
#1;data_in = testData4[950];
@(posedge clk);
#1;data_in = testData4[951];
@(posedge clk);
#1;data_in = testData4[952];
@(posedge clk);
#1;data_in = testData4[953];
@(posedge clk);
#1;data_in = testData4[954];
@(posedge clk);
#1;data_in = testData4[955];
@(posedge clk);
#1;data_in = testData4[956];
@(posedge clk);
#1;data_in = testData4[957];
@(posedge clk);
#1;data_in = testData4[958];
@(posedge clk);
#1;data_in = testData4[959];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[960]; 
@(posedge clk);
#1;data_in = testData4[961];
@(posedge clk);
#1;data_in = testData4[962];
@(posedge clk);
#1;data_in = testData4[963];
@(posedge clk);
#1;data_in = testData4[964];
@(posedge clk);
#1;data_in = testData4[965];
@(posedge clk);
#1;data_in = testData4[966];
@(posedge clk);
#1;data_in = testData4[967];
@(posedge clk);
#1;data_in = testData4[968];
@(posedge clk);
#1;data_in = testData4[969];
@(posedge clk);
#1;data_in = testData4[970];
@(posedge clk);
#1;data_in = testData4[971];
@(posedge clk);
#1;data_in = testData4[972];
@(posedge clk);
#1;data_in = testData4[973];
@(posedge clk);
#1;data_in = testData4[974];
@(posedge clk);
#1;data_in = testData4[975];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[976]; 
@(posedge clk);
#1;data_in = testData4[977];
@(posedge clk);
#1;data_in = testData4[978];
@(posedge clk);
#1;data_in = testData4[979];
@(posedge clk);
#1;data_in = testData4[980];
@(posedge clk);
#1;data_in = testData4[981];
@(posedge clk);
#1;data_in = testData4[982];
@(posedge clk);
#1;data_in = testData4[983];
@(posedge clk);
#1;data_in = testData4[984];
@(posedge clk);
#1;data_in = testData4[985];
@(posedge clk);
#1;data_in = testData4[986];
@(posedge clk);
#1;data_in = testData4[987];
@(posedge clk);
#1;data_in = testData4[988];
@(posedge clk);
#1;data_in = testData4[989];
@(posedge clk);
#1;data_in = testData4[990];
@(posedge clk);
#1;data_in = testData4[991];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[992]; 
@(posedge clk);
#1;data_in = testData4[993];
@(posedge clk);
#1;data_in = testData4[994];
@(posedge clk);
#1;data_in = testData4[995];
@(posedge clk);
#1;data_in = testData4[996];
@(posedge clk);
#1;data_in = testData4[997];
@(posedge clk);
#1;data_in = testData4[998];
@(posedge clk);
#1;data_in = testData4[999];
@(posedge clk);
#1;data_in = testData4[1000];
@(posedge clk);
#1;data_in = testData4[1001];
@(posedge clk);
#1;data_in = testData4[1002];
@(posedge clk);
#1;data_in = testData4[1003];
@(posedge clk);
#1;data_in = testData4[1004];
@(posedge clk);
#1;data_in = testData4[1005];
@(posedge clk);
#1;data_in = testData4[1006];
@(posedge clk);
#1;data_in = testData4[1007];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[1008]; 
@(posedge clk);
#1;data_in = testData4[1009];
@(posedge clk);
#1;data_in = testData4[1010];
@(posedge clk);
#1;data_in = testData4[1011];
@(posedge clk);
#1;data_in = testData4[1012];
@(posedge clk);
#1;data_in = testData4[1013];
@(posedge clk);
#1;data_in = testData4[1014];
@(posedge clk);
#1;data_in = testData4[1015];
@(posedge clk);
#1;data_in = testData4[1016];
@(posedge clk);
#1;data_in = testData4[1017];
@(posedge clk);
#1;data_in = testData4[1018];
@(posedge clk);
#1;data_in = testData4[1019];
@(posedge clk);
#1;data_in = testData4[1020];
@(posedge clk);
#1;data_in = testData4[1021];
@(posedge clk);
#1;data_in = testData4[1022];
@(posedge clk);
#1;data_in = testData4[1023];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[1024]; 
@(posedge clk);
#1;data_in = testData4[1025];
@(posedge clk);
#1;data_in = testData4[1026];
@(posedge clk);
#1;data_in = testData4[1027];
@(posedge clk);
#1;data_in = testData4[1028];
@(posedge clk);
#1;data_in = testData4[1029];
@(posedge clk);
#1;data_in = testData4[1030];
@(posedge clk);
#1;data_in = testData4[1031];
@(posedge clk);
#1;data_in = testData4[1032];
@(posedge clk);
#1;data_in = testData4[1033];
@(posedge clk);
#1;data_in = testData4[1034];
@(posedge clk);
#1;data_in = testData4[1035];
@(posedge clk);
#1;data_in = testData4[1036];
@(posedge clk);
#1;data_in = testData4[1037];
@(posedge clk);
#1;data_in = testData4[1038];
@(posedge clk);
#1;data_in = testData4[1039];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[1040]; 
@(posedge clk);
#1;data_in = testData4[1041];
@(posedge clk);
#1;data_in = testData4[1042];
@(posedge clk);
#1;data_in = testData4[1043];
@(posedge clk);
#1;data_in = testData4[1044];
@(posedge clk);
#1;data_in = testData4[1045];
@(posedge clk);
#1;data_in = testData4[1046];
@(posedge clk);
#1;data_in = testData4[1047];
@(posedge clk);
#1;data_in = testData4[1048];
@(posedge clk);
#1;data_in = testData4[1049];
@(posedge clk);
#1;data_in = testData4[1050];
@(posedge clk);
#1;data_in = testData4[1051];
@(posedge clk);
#1;data_in = testData4[1052];
@(posedge clk);
#1;data_in = testData4[1053];
@(posedge clk);
#1;data_in = testData4[1054];
@(posedge clk);
#1;data_in = testData4[1055];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[1056]; 
@(posedge clk);
#1;data_in = testData4[1057];
@(posedge clk);
#1;data_in = testData4[1058];
@(posedge clk);
#1;data_in = testData4[1059];
@(posedge clk);
#1;data_in = testData4[1060];
@(posedge clk);
#1;data_in = testData4[1061];
@(posedge clk);
#1;data_in = testData4[1062];
@(posedge clk);
#1;data_in = testData4[1063];
@(posedge clk);
#1;data_in = testData4[1064];
@(posedge clk);
#1;data_in = testData4[1065];
@(posedge clk);
#1;data_in = testData4[1066];
@(posedge clk);
#1;data_in = testData4[1067];
@(posedge clk);
#1;data_in = testData4[1068];
@(posedge clk);
#1;data_in = testData4[1069];
@(posedge clk);
#1;data_in = testData4[1070];
@(posedge clk);
#1;data_in = testData4[1071];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
module tb6();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData6[13871:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb6", testData6);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb6");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[0];
@(posedge clk);
#1;data_in = testData6[1];
@(posedge clk);
#1;data_in = testData6[2];
@(posedge clk);
#1;data_in = testData6[3];
@(posedge clk);
#1;data_in = testData6[4];
@(posedge clk);
#1;data_in = testData6[5];
@(posedge clk);
#1;data_in = testData6[6];
@(posedge clk);
#1;data_in = testData6[7];
@(posedge clk);
#1;data_in = testData6[8];
@(posedge clk);
#1;data_in = testData6[9];
@(posedge clk);
#1;data_in = testData6[10];
@(posedge clk);
#1;data_in = testData6[11];
@(posedge clk);
#1;data_in = testData6[12];
@(posedge clk);
#1;data_in = testData6[13];
@(posedge clk);
#1;data_in = testData6[14];
@(posedge clk);
#1;data_in = testData6[15];
@(posedge clk);
#1;data_in = testData6[16];
@(posedge clk);
#1;data_in = testData6[17];
@(posedge clk);
#1;data_in = testData6[18];
@(posedge clk);
#1;data_in = testData6[19];
@(posedge clk);
#1;data_in = testData6[20];
@(posedge clk);
#1;data_in = testData6[21];
@(posedge clk);
#1;data_in = testData6[22];
@(posedge clk);
#1;data_in = testData6[23];
@(posedge clk);
#1;data_in = testData6[24];
@(posedge clk);
#1;data_in = testData6[25];
@(posedge clk);
#1;data_in = testData6[26];
@(posedge clk);
#1;data_in = testData6[27];
@(posedge clk);
#1;data_in = testData6[28];
@(posedge clk);
#1;data_in = testData6[29];
@(posedge clk);
#1;data_in = testData6[30];
@(posedge clk);
#1;data_in = testData6[31];
@(posedge clk);
#1;data_in = testData6[32];
@(posedge clk);
#1;data_in = testData6[33];
@(posedge clk);
#1;data_in = testData6[34];
@(posedge clk);
#1;data_in = testData6[35];
@(posedge clk);
#1;data_in = testData6[36];
@(posedge clk);
#1;data_in = testData6[37];
@(posedge clk);
#1;data_in = testData6[38];
@(posedge clk);
#1;data_in = testData6[39];
@(posedge clk);
#1;data_in = testData6[40];
@(posedge clk);
#1;data_in = testData6[41];
@(posedge clk);
#1;data_in = testData6[42];
@(posedge clk);
#1;data_in = testData6[43];
@(posedge clk);
#1;data_in = testData6[44];
@(posedge clk);
#1;data_in = testData6[45];
@(posedge clk);
#1;data_in = testData6[46];
@(posedge clk);
#1;data_in = testData6[47];
@(posedge clk);
#1;data_in = testData6[48];
@(posedge clk);
#1;data_in = testData6[49];
@(posedge clk);
#1;data_in = testData6[50];
@(posedge clk);
#1;data_in = testData6[51];
@(posedge clk);
#1;data_in = testData6[52];
@(posedge clk);
#1;data_in = testData6[53];
@(posedge clk);
#1;data_in = testData6[54];
@(posedge clk);
#1;data_in = testData6[55];
@(posedge clk);
#1;data_in = testData6[56];
@(posedge clk);
#1;data_in = testData6[57];
@(posedge clk);
#1;data_in = testData6[58];
@(posedge clk);
#1;data_in = testData6[59];
@(posedge clk);
#1;data_in = testData6[60];
@(posedge clk);
#1;data_in = testData6[61];
@(posedge clk);
#1;data_in = testData6[62];
@(posedge clk);
#1;data_in = testData6[63];
@(posedge clk);
#1;data_in = testData6[64];
@(posedge clk);
#1;data_in = testData6[65];
@(posedge clk);
#1;data_in = testData6[66];
@(posedge clk);
#1;data_in = testData6[67];
@(posedge clk);
#1;data_in = testData6[68];
@(posedge clk);
#1;data_in = testData6[69];
@(posedge clk);
#1;data_in = testData6[70];
@(posedge clk);
#1;data_in = testData6[71];
@(posedge clk);
#1;data_in = testData6[72];
@(posedge clk);
#1;data_in = testData6[73];
@(posedge clk);
#1;data_in = testData6[74];
@(posedge clk);
#1;data_in = testData6[75];
@(posedge clk);
#1;data_in = testData6[76];
@(posedge clk);
#1;data_in = testData6[77];
@(posedge clk);
#1;data_in = testData6[78];
@(posedge clk);
#1;data_in = testData6[79];
@(posedge clk);
#1;data_in = testData6[80];
@(posedge clk);
#1;data_in = testData6[81];
@(posedge clk);
#1;data_in = testData6[82];
@(posedge clk);
#1;data_in = testData6[83];
@(posedge clk);
#1;data_in = testData6[84];
@(posedge clk);
#1;data_in = testData6[85];
@(posedge clk);
#1;data_in = testData6[86];
@(posedge clk);
#1;data_in = testData6[87];
@(posedge clk);
#1;data_in = testData6[88];
@(posedge clk);
#1;data_in = testData6[89];
@(posedge clk);
#1;data_in = testData6[90];
@(posedge clk);
#1;data_in = testData6[91];
@(posedge clk);
#1;data_in = testData6[92];
@(posedge clk);
#1;data_in = testData6[93];
@(posedge clk);
#1;data_in = testData6[94];
@(posedge clk);
#1;data_in = testData6[95];
@(posedge clk);
#1;data_in = testData6[96];
@(posedge clk);
#1;data_in = testData6[97];
@(posedge clk);
#1;data_in = testData6[98];
@(posedge clk);
#1;data_in = testData6[99];
@(posedge clk);
#1;data_in = testData6[100];
@(posedge clk);
#1;data_in = testData6[101];
@(posedge clk);
#1;data_in = testData6[102];
@(posedge clk);
#1;data_in = testData6[103];
@(posedge clk);
#1;data_in = testData6[104];
@(posedge clk);
#1;data_in = testData6[105];
@(posedge clk);
#1;data_in = testData6[106];
@(posedge clk);
#1;data_in = testData6[107];
@(posedge clk);
#1;data_in = testData6[108];
@(posedge clk);
#1;data_in = testData6[109];
@(posedge clk);
#1;data_in = testData6[110];
@(posedge clk);
#1;data_in = testData6[111];
@(posedge clk);
#1;data_in = testData6[112];
@(posedge clk);
#1;data_in = testData6[113];
@(posedge clk);
#1;data_in = testData6[114];
@(posedge clk);
#1;data_in = testData6[115];
@(posedge clk);
#1;data_in = testData6[116];
@(posedge clk);
#1;data_in = testData6[117];
@(posedge clk);
#1;data_in = testData6[118];
@(posedge clk);
#1;data_in = testData6[119];
@(posedge clk);
#1;data_in = testData6[120];
@(posedge clk);
#1;data_in = testData6[121];
@(posedge clk);
#1;data_in = testData6[122];
@(posedge clk);
#1;data_in = testData6[123];
@(posedge clk);
#1;data_in = testData6[124];
@(posedge clk);
#1;data_in = testData6[125];
@(posedge clk);
#1;data_in = testData6[126];
@(posedge clk);
#1;data_in = testData6[127];
@(posedge clk);
#1;data_in = testData6[128];
@(posedge clk);
#1;data_in = testData6[129];
@(posedge clk);
#1;data_in = testData6[130];
@(posedge clk);
#1;data_in = testData6[131];
@(posedge clk);
#1;data_in = testData6[132];
@(posedge clk);
#1;data_in = testData6[133];
@(posedge clk);
#1;data_in = testData6[134];
@(posedge clk);
#1;data_in = testData6[135];
@(posedge clk);
#1;data_in = testData6[136];
@(posedge clk);
#1;data_in = testData6[137];
@(posedge clk);
#1;data_in = testData6[138];
@(posedge clk);
#1;data_in = testData6[139];
@(posedge clk);
#1;data_in = testData6[140];
@(posedge clk);
#1;data_in = testData6[141];
@(posedge clk);
#1;data_in = testData6[142];
@(posedge clk);
#1;data_in = testData6[143];
@(posedge clk);
#1;data_in = testData6[144];
@(posedge clk);
#1;data_in = testData6[145];
@(posedge clk);
#1;data_in = testData6[146];
@(posedge clk);
#1;data_in = testData6[147];
@(posedge clk);
#1;data_in = testData6[148];
@(posedge clk);
#1;data_in = testData6[149];
@(posedge clk);
#1;data_in = testData6[150];
@(posedge clk);
#1;data_in = testData6[151];
@(posedge clk);
#1;data_in = testData6[152];
@(posedge clk);
#1;data_in = testData6[153];
@(posedge clk);
#1;data_in = testData6[154];
@(posedge clk);
#1;data_in = testData6[155];
@(posedge clk);
#1;data_in = testData6[156];
@(posedge clk);
#1;data_in = testData6[157];
@(posedge clk);
#1;data_in = testData6[158];
@(posedge clk);
#1;data_in = testData6[159];
@(posedge clk);
#1;data_in = testData6[160];
@(posedge clk);
#1;data_in = testData6[161];
@(posedge clk);
#1;data_in = testData6[162];
@(posedge clk);
#1;data_in = testData6[163];
@(posedge clk);
#1;data_in = testData6[164];
@(posedge clk);
#1;data_in = testData6[165];
@(posedge clk);
#1;data_in = testData6[166];
@(posedge clk);
#1;data_in = testData6[167];
@(posedge clk);
#1;data_in = testData6[168];
@(posedge clk);
#1;data_in = testData6[169];
@(posedge clk);
#1;data_in = testData6[170];
@(posedge clk);
#1;data_in = testData6[171];
@(posedge clk);
#1;data_in = testData6[172];
@(posedge clk);
#1;data_in = testData6[173];
@(posedge clk);
#1;data_in = testData6[174];
@(posedge clk);
#1;data_in = testData6[175];
@(posedge clk);
#1;data_in = testData6[176];
@(posedge clk);
#1;data_in = testData6[177];
@(posedge clk);
#1;data_in = testData6[178];
@(posedge clk);
#1;data_in = testData6[179];
@(posedge clk);
#1;data_in = testData6[180];
@(posedge clk);
#1;data_in = testData6[181];
@(posedge clk);
#1;data_in = testData6[182];
@(posedge clk);
#1;data_in = testData6[183];
@(posedge clk);
#1;data_in = testData6[184];
@(posedge clk);
#1;data_in = testData6[185];
@(posedge clk);
#1;data_in = testData6[186];
@(posedge clk);
#1;data_in = testData6[187];
@(posedge clk);
#1;data_in = testData6[188];
@(posedge clk);
#1;data_in = testData6[189];
@(posedge clk);
#1;data_in = testData6[190];
@(posedge clk);
#1;data_in = testData6[191];
@(posedge clk);
#1;data_in = testData6[192];
@(posedge clk);
#1;data_in = testData6[193];
@(posedge clk);
#1;data_in = testData6[194];
@(posedge clk);
#1;data_in = testData6[195];
@(posedge clk);
#1;data_in = testData6[196];
@(posedge clk);
#1;data_in = testData6[197];
@(posedge clk);
#1;data_in = testData6[198];
@(posedge clk);
#1;data_in = testData6[199];
@(posedge clk);
#1;data_in = testData6[200];
@(posedge clk);
#1;data_in = testData6[201];
@(posedge clk);
#1;data_in = testData6[202];
@(posedge clk);
#1;data_in = testData6[203];
@(posedge clk);
#1;data_in = testData6[204];
@(posedge clk);
#1;data_in = testData6[205];
@(posedge clk);
#1;data_in = testData6[206];
@(posedge clk);
#1;data_in = testData6[207];
@(posedge clk);
#1;data_in = testData6[208];
@(posedge clk);
#1;data_in = testData6[209];
@(posedge clk);
#1;data_in = testData6[210];
@(posedge clk);
#1;data_in = testData6[211];
@(posedge clk);
#1;data_in = testData6[212];
@(posedge clk);
#1;data_in = testData6[213];
@(posedge clk);
#1;data_in = testData6[214];
@(posedge clk);
#1;data_in = testData6[215];
@(posedge clk);
#1;data_in = testData6[216];
@(posedge clk);
#1;data_in = testData6[217];
@(posedge clk);
#1;data_in = testData6[218];
@(posedge clk);
#1;data_in = testData6[219];
@(posedge clk);
#1;data_in = testData6[220];
@(posedge clk);
#1;data_in = testData6[221];
@(posedge clk);
#1;data_in = testData6[222];
@(posedge clk);
#1;data_in = testData6[223];
@(posedge clk);
#1;data_in = testData6[224];
@(posedge clk);
#1;data_in = testData6[225];
@(posedge clk);
#1;data_in = testData6[226];
@(posedge clk);
#1;data_in = testData6[227];
@(posedge clk);
#1;data_in = testData6[228];
@(posedge clk);
#1;data_in = testData6[229];
@(posedge clk);
#1;data_in = testData6[230];
@(posedge clk);
#1;data_in = testData6[231];
@(posedge clk);
#1;data_in = testData6[232];
@(posedge clk);
#1;data_in = testData6[233];
@(posedge clk);
#1;data_in = testData6[234];
@(posedge clk);
#1;data_in = testData6[235];
@(posedge clk);
#1;data_in = testData6[236];
@(posedge clk);
#1;data_in = testData6[237];
@(posedge clk);
#1;data_in = testData6[238];
@(posedge clk);
#1;data_in = testData6[239];
@(posedge clk);
#1;data_in = testData6[240];
@(posedge clk);
#1;data_in = testData6[241];
@(posedge clk);
#1;data_in = testData6[242];
@(posedge clk);
#1;data_in = testData6[243];
@(posedge clk);
#1;data_in = testData6[244];
@(posedge clk);
#1;data_in = testData6[245];
@(posedge clk);
#1;data_in = testData6[246];
@(posedge clk);
#1;data_in = testData6[247];
@(posedge clk);
#1;data_in = testData6[248];
@(posedge clk);
#1;data_in = testData6[249];
@(posedge clk);
#1;data_in = testData6[250];
@(posedge clk);
#1;data_in = testData6[251];
@(posedge clk);
#1;data_in = testData6[252];
@(posedge clk);
#1;data_in = testData6[253];
@(posedge clk);
#1;data_in = testData6[254];
@(posedge clk);
#1;data_in = testData6[255];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[256]; 
@(posedge clk);
#1;data_in = testData6[257];
@(posedge clk);
#1;data_in = testData6[258];
@(posedge clk);
#1;data_in = testData6[259];
@(posedge clk);
#1;data_in = testData6[260];
@(posedge clk);
#1;data_in = testData6[261];
@(posedge clk);
#1;data_in = testData6[262];
@(posedge clk);
#1;data_in = testData6[263];
@(posedge clk);
#1;data_in = testData6[264];
@(posedge clk);
#1;data_in = testData6[265];
@(posedge clk);
#1;data_in = testData6[266];
@(posedge clk);
#1;data_in = testData6[267];
@(posedge clk);
#1;data_in = testData6[268];
@(posedge clk);
#1;data_in = testData6[269];
@(posedge clk);
#1;data_in = testData6[270];
@(posedge clk);
#1;data_in = testData6[271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[272];
@(posedge clk);
#1;data_in = testData6[273];
@(posedge clk);
#1;data_in = testData6[274];
@(posedge clk);
#1;data_in = testData6[275];
@(posedge clk);
#1;data_in = testData6[276];
@(posedge clk);
#1;data_in = testData6[277];
@(posedge clk);
#1;data_in = testData6[278];
@(posedge clk);
#1;data_in = testData6[279];
@(posedge clk);
#1;data_in = testData6[280];
@(posedge clk);
#1;data_in = testData6[281];
@(posedge clk);
#1;data_in = testData6[282];
@(posedge clk);
#1;data_in = testData6[283];
@(posedge clk);
#1;data_in = testData6[284];
@(posedge clk);
#1;data_in = testData6[285];
@(posedge clk);
#1;data_in = testData6[286];
@(posedge clk);
#1;data_in = testData6[287];
@(posedge clk);
#1;data_in = testData6[288];
@(posedge clk);
#1;data_in = testData6[289];
@(posedge clk);
#1;data_in = testData6[290];
@(posedge clk);
#1;data_in = testData6[291];
@(posedge clk);
#1;data_in = testData6[292];
@(posedge clk);
#1;data_in = testData6[293];
@(posedge clk);
#1;data_in = testData6[294];
@(posedge clk);
#1;data_in = testData6[295];
@(posedge clk);
#1;data_in = testData6[296];
@(posedge clk);
#1;data_in = testData6[297];
@(posedge clk);
#1;data_in = testData6[298];
@(posedge clk);
#1;data_in = testData6[299];
@(posedge clk);
#1;data_in = testData6[300];
@(posedge clk);
#1;data_in = testData6[301];
@(posedge clk);
#1;data_in = testData6[302];
@(posedge clk);
#1;data_in = testData6[303];
@(posedge clk);
#1;data_in = testData6[304];
@(posedge clk);
#1;data_in = testData6[305];
@(posedge clk);
#1;data_in = testData6[306];
@(posedge clk);
#1;data_in = testData6[307];
@(posedge clk);
#1;data_in = testData6[308];
@(posedge clk);
#1;data_in = testData6[309];
@(posedge clk);
#1;data_in = testData6[310];
@(posedge clk);
#1;data_in = testData6[311];
@(posedge clk);
#1;data_in = testData6[312];
@(posedge clk);
#1;data_in = testData6[313];
@(posedge clk);
#1;data_in = testData6[314];
@(posedge clk);
#1;data_in = testData6[315];
@(posedge clk);
#1;data_in = testData6[316];
@(posedge clk);
#1;data_in = testData6[317];
@(posedge clk);
#1;data_in = testData6[318];
@(posedge clk);
#1;data_in = testData6[319];
@(posedge clk);
#1;data_in = testData6[320];
@(posedge clk);
#1;data_in = testData6[321];
@(posedge clk);
#1;data_in = testData6[322];
@(posedge clk);
#1;data_in = testData6[323];
@(posedge clk);
#1;data_in = testData6[324];
@(posedge clk);
#1;data_in = testData6[325];
@(posedge clk);
#1;data_in = testData6[326];
@(posedge clk);
#1;data_in = testData6[327];
@(posedge clk);
#1;data_in = testData6[328];
@(posedge clk);
#1;data_in = testData6[329];
@(posedge clk);
#1;data_in = testData6[330];
@(posedge clk);
#1;data_in = testData6[331];
@(posedge clk);
#1;data_in = testData6[332];
@(posedge clk);
#1;data_in = testData6[333];
@(posedge clk);
#1;data_in = testData6[334];
@(posedge clk);
#1;data_in = testData6[335];
@(posedge clk);
#1;data_in = testData6[336];
@(posedge clk);
#1;data_in = testData6[337];
@(posedge clk);
#1;data_in = testData6[338];
@(posedge clk);
#1;data_in = testData6[339];
@(posedge clk);
#1;data_in = testData6[340];
@(posedge clk);
#1;data_in = testData6[341];
@(posedge clk);
#1;data_in = testData6[342];
@(posedge clk);
#1;data_in = testData6[343];
@(posedge clk);
#1;data_in = testData6[344];
@(posedge clk);
#1;data_in = testData6[345];
@(posedge clk);
#1;data_in = testData6[346];
@(posedge clk);
#1;data_in = testData6[347];
@(posedge clk);
#1;data_in = testData6[348];
@(posedge clk);
#1;data_in = testData6[349];
@(posedge clk);
#1;data_in = testData6[350];
@(posedge clk);
#1;data_in = testData6[351];
@(posedge clk);
#1;data_in = testData6[352];
@(posedge clk);
#1;data_in = testData6[353];
@(posedge clk);
#1;data_in = testData6[354];
@(posedge clk);
#1;data_in = testData6[355];
@(posedge clk);
#1;data_in = testData6[356];
@(posedge clk);
#1;data_in = testData6[357];
@(posedge clk);
#1;data_in = testData6[358];
@(posedge clk);
#1;data_in = testData6[359];
@(posedge clk);
#1;data_in = testData6[360];
@(posedge clk);
#1;data_in = testData6[361];
@(posedge clk);
#1;data_in = testData6[362];
@(posedge clk);
#1;data_in = testData6[363];
@(posedge clk);
#1;data_in = testData6[364];
@(posedge clk);
#1;data_in = testData6[365];
@(posedge clk);
#1;data_in = testData6[366];
@(posedge clk);
#1;data_in = testData6[367];
@(posedge clk);
#1;data_in = testData6[368];
@(posedge clk);
#1;data_in = testData6[369];
@(posedge clk);
#1;data_in = testData6[370];
@(posedge clk);
#1;data_in = testData6[371];
@(posedge clk);
#1;data_in = testData6[372];
@(posedge clk);
#1;data_in = testData6[373];
@(posedge clk);
#1;data_in = testData6[374];
@(posedge clk);
#1;data_in = testData6[375];
@(posedge clk);
#1;data_in = testData6[376];
@(posedge clk);
#1;data_in = testData6[377];
@(posedge clk);
#1;data_in = testData6[378];
@(posedge clk);
#1;data_in = testData6[379];
@(posedge clk);
#1;data_in = testData6[380];
@(posedge clk);
#1;data_in = testData6[381];
@(posedge clk);
#1;data_in = testData6[382];
@(posedge clk);
#1;data_in = testData6[383];
@(posedge clk);
#1;data_in = testData6[384];
@(posedge clk);
#1;data_in = testData6[385];
@(posedge clk);
#1;data_in = testData6[386];
@(posedge clk);
#1;data_in = testData6[387];
@(posedge clk);
#1;data_in = testData6[388];
@(posedge clk);
#1;data_in = testData6[389];
@(posedge clk);
#1;data_in = testData6[390];
@(posedge clk);
#1;data_in = testData6[391];
@(posedge clk);
#1;data_in = testData6[392];
@(posedge clk);
#1;data_in = testData6[393];
@(posedge clk);
#1;data_in = testData6[394];
@(posedge clk);
#1;data_in = testData6[395];
@(posedge clk);
#1;data_in = testData6[396];
@(posedge clk);
#1;data_in = testData6[397];
@(posedge clk);
#1;data_in = testData6[398];
@(posedge clk);
#1;data_in = testData6[399];
@(posedge clk);
#1;data_in = testData6[400];
@(posedge clk);
#1;data_in = testData6[401];
@(posedge clk);
#1;data_in = testData6[402];
@(posedge clk);
#1;data_in = testData6[403];
@(posedge clk);
#1;data_in = testData6[404];
@(posedge clk);
#1;data_in = testData6[405];
@(posedge clk);
#1;data_in = testData6[406];
@(posedge clk);
#1;data_in = testData6[407];
@(posedge clk);
#1;data_in = testData6[408];
@(posedge clk);
#1;data_in = testData6[409];
@(posedge clk);
#1;data_in = testData6[410];
@(posedge clk);
#1;data_in = testData6[411];
@(posedge clk);
#1;data_in = testData6[412];
@(posedge clk);
#1;data_in = testData6[413];
@(posedge clk);
#1;data_in = testData6[414];
@(posedge clk);
#1;data_in = testData6[415];
@(posedge clk);
#1;data_in = testData6[416];
@(posedge clk);
#1;data_in = testData6[417];
@(posedge clk);
#1;data_in = testData6[418];
@(posedge clk);
#1;data_in = testData6[419];
@(posedge clk);
#1;data_in = testData6[420];
@(posedge clk);
#1;data_in = testData6[421];
@(posedge clk);
#1;data_in = testData6[422];
@(posedge clk);
#1;data_in = testData6[423];
@(posedge clk);
#1;data_in = testData6[424];
@(posedge clk);
#1;data_in = testData6[425];
@(posedge clk);
#1;data_in = testData6[426];
@(posedge clk);
#1;data_in = testData6[427];
@(posedge clk);
#1;data_in = testData6[428];
@(posedge clk);
#1;data_in = testData6[429];
@(posedge clk);
#1;data_in = testData6[430];
@(posedge clk);
#1;data_in = testData6[431];
@(posedge clk);
#1;data_in = testData6[432];
@(posedge clk);
#1;data_in = testData6[433];
@(posedge clk);
#1;data_in = testData6[434];
@(posedge clk);
#1;data_in = testData6[435];
@(posedge clk);
#1;data_in = testData6[436];
@(posedge clk);
#1;data_in = testData6[437];
@(posedge clk);
#1;data_in = testData6[438];
@(posedge clk);
#1;data_in = testData6[439];
@(posedge clk);
#1;data_in = testData6[440];
@(posedge clk);
#1;data_in = testData6[441];
@(posedge clk);
#1;data_in = testData6[442];
@(posedge clk);
#1;data_in = testData6[443];
@(posedge clk);
#1;data_in = testData6[444];
@(posedge clk);
#1;data_in = testData6[445];
@(posedge clk);
#1;data_in = testData6[446];
@(posedge clk);
#1;data_in = testData6[447];
@(posedge clk);
#1;data_in = testData6[448];
@(posedge clk);
#1;data_in = testData6[449];
@(posedge clk);
#1;data_in = testData6[450];
@(posedge clk);
#1;data_in = testData6[451];
@(posedge clk);
#1;data_in = testData6[452];
@(posedge clk);
#1;data_in = testData6[453];
@(posedge clk);
#1;data_in = testData6[454];
@(posedge clk);
#1;data_in = testData6[455];
@(posedge clk);
#1;data_in = testData6[456];
@(posedge clk);
#1;data_in = testData6[457];
@(posedge clk);
#1;data_in = testData6[458];
@(posedge clk);
#1;data_in = testData6[459];
@(posedge clk);
#1;data_in = testData6[460];
@(posedge clk);
#1;data_in = testData6[461];
@(posedge clk);
#1;data_in = testData6[462];
@(posedge clk);
#1;data_in = testData6[463];
@(posedge clk);
#1;data_in = testData6[464];
@(posedge clk);
#1;data_in = testData6[465];
@(posedge clk);
#1;data_in = testData6[466];
@(posedge clk);
#1;data_in = testData6[467];
@(posedge clk);
#1;data_in = testData6[468];
@(posedge clk);
#1;data_in = testData6[469];
@(posedge clk);
#1;data_in = testData6[470];
@(posedge clk);
#1;data_in = testData6[471];
@(posedge clk);
#1;data_in = testData6[472];
@(posedge clk);
#1;data_in = testData6[473];
@(posedge clk);
#1;data_in = testData6[474];
@(posedge clk);
#1;data_in = testData6[475];
@(posedge clk);
#1;data_in = testData6[476];
@(posedge clk);
#1;data_in = testData6[477];
@(posedge clk);
#1;data_in = testData6[478];
@(posedge clk);
#1;data_in = testData6[479];
@(posedge clk);
#1;data_in = testData6[480];
@(posedge clk);
#1;data_in = testData6[481];
@(posedge clk);
#1;data_in = testData6[482];
@(posedge clk);
#1;data_in = testData6[483];
@(posedge clk);
#1;data_in = testData6[484];
@(posedge clk);
#1;data_in = testData6[485];
@(posedge clk);
#1;data_in = testData6[486];
@(posedge clk);
#1;data_in = testData6[487];
@(posedge clk);
#1;data_in = testData6[488];
@(posedge clk);
#1;data_in = testData6[489];
@(posedge clk);
#1;data_in = testData6[490];
@(posedge clk);
#1;data_in = testData6[491];
@(posedge clk);
#1;data_in = testData6[492];
@(posedge clk);
#1;data_in = testData6[493];
@(posedge clk);
#1;data_in = testData6[494];
@(posedge clk);
#1;data_in = testData6[495];
@(posedge clk);
#1;data_in = testData6[496];
@(posedge clk);
#1;data_in = testData6[497];
@(posedge clk);
#1;data_in = testData6[498];
@(posedge clk);
#1;data_in = testData6[499];
@(posedge clk);
#1;data_in = testData6[500];
@(posedge clk);
#1;data_in = testData6[501];
@(posedge clk);
#1;data_in = testData6[502];
@(posedge clk);
#1;data_in = testData6[503];
@(posedge clk);
#1;data_in = testData6[504];
@(posedge clk);
#1;data_in = testData6[505];
@(posedge clk);
#1;data_in = testData6[506];
@(posedge clk);
#1;data_in = testData6[507];
@(posedge clk);
#1;data_in = testData6[508];
@(posedge clk);
#1;data_in = testData6[509];
@(posedge clk);
#1;data_in = testData6[510];
@(posedge clk);
#1;data_in = testData6[511];
@(posedge clk);
#1;data_in = testData6[512];
@(posedge clk);
#1;data_in = testData6[513];
@(posedge clk);
#1;data_in = testData6[514];
@(posedge clk);
#1;data_in = testData6[515];
@(posedge clk);
#1;data_in = testData6[516];
@(posedge clk);
#1;data_in = testData6[517];
@(posedge clk);
#1;data_in = testData6[518];
@(posedge clk);
#1;data_in = testData6[519];
@(posedge clk);
#1;data_in = testData6[520];
@(posedge clk);
#1;data_in = testData6[521];
@(posedge clk);
#1;data_in = testData6[522];
@(posedge clk);
#1;data_in = testData6[523];
@(posedge clk);
#1;data_in = testData6[524];
@(posedge clk);
#1;data_in = testData6[525];
@(posedge clk);
#1;data_in = testData6[526];
@(posedge clk);
#1;data_in = testData6[527];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[528]; 
@(posedge clk);
#1;data_in = testData6[529];
@(posedge clk);
#1;data_in = testData6[530];
@(posedge clk);
#1;data_in = testData6[531];
@(posedge clk);
#1;data_in = testData6[532];
@(posedge clk);
#1;data_in = testData6[533];
@(posedge clk);
#1;data_in = testData6[534];
@(posedge clk);
#1;data_in = testData6[535];
@(posedge clk);
#1;data_in = testData6[536];
@(posedge clk);
#1;data_in = testData6[537];
@(posedge clk);
#1;data_in = testData6[538];
@(posedge clk);
#1;data_in = testData6[539];
@(posedge clk);
#1;data_in = testData6[540];
@(posedge clk);
#1;data_in = testData6[541];
@(posedge clk);
#1;data_in = testData6[542];
@(posedge clk);
#1;data_in = testData6[543];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[544];
@(posedge clk);
#1;data_in = testData6[545];
@(posedge clk);
#1;data_in = testData6[546];
@(posedge clk);
#1;data_in = testData6[547];
@(posedge clk);
#1;data_in = testData6[548];
@(posedge clk);
#1;data_in = testData6[549];
@(posedge clk);
#1;data_in = testData6[550];
@(posedge clk);
#1;data_in = testData6[551];
@(posedge clk);
#1;data_in = testData6[552];
@(posedge clk);
#1;data_in = testData6[553];
@(posedge clk);
#1;data_in = testData6[554];
@(posedge clk);
#1;data_in = testData6[555];
@(posedge clk);
#1;data_in = testData6[556];
@(posedge clk);
#1;data_in = testData6[557];
@(posedge clk);
#1;data_in = testData6[558];
@(posedge clk);
#1;data_in = testData6[559];
@(posedge clk);
#1;data_in = testData6[560];
@(posedge clk);
#1;data_in = testData6[561];
@(posedge clk);
#1;data_in = testData6[562];
@(posedge clk);
#1;data_in = testData6[563];
@(posedge clk);
#1;data_in = testData6[564];
@(posedge clk);
#1;data_in = testData6[565];
@(posedge clk);
#1;data_in = testData6[566];
@(posedge clk);
#1;data_in = testData6[567];
@(posedge clk);
#1;data_in = testData6[568];
@(posedge clk);
#1;data_in = testData6[569];
@(posedge clk);
#1;data_in = testData6[570];
@(posedge clk);
#1;data_in = testData6[571];
@(posedge clk);
#1;data_in = testData6[572];
@(posedge clk);
#1;data_in = testData6[573];
@(posedge clk);
#1;data_in = testData6[574];
@(posedge clk);
#1;data_in = testData6[575];
@(posedge clk);
#1;data_in = testData6[576];
@(posedge clk);
#1;data_in = testData6[577];
@(posedge clk);
#1;data_in = testData6[578];
@(posedge clk);
#1;data_in = testData6[579];
@(posedge clk);
#1;data_in = testData6[580];
@(posedge clk);
#1;data_in = testData6[581];
@(posedge clk);
#1;data_in = testData6[582];
@(posedge clk);
#1;data_in = testData6[583];
@(posedge clk);
#1;data_in = testData6[584];
@(posedge clk);
#1;data_in = testData6[585];
@(posedge clk);
#1;data_in = testData6[586];
@(posedge clk);
#1;data_in = testData6[587];
@(posedge clk);
#1;data_in = testData6[588];
@(posedge clk);
#1;data_in = testData6[589];
@(posedge clk);
#1;data_in = testData6[590];
@(posedge clk);
#1;data_in = testData6[591];
@(posedge clk);
#1;data_in = testData6[592];
@(posedge clk);
#1;data_in = testData6[593];
@(posedge clk);
#1;data_in = testData6[594];
@(posedge clk);
#1;data_in = testData6[595];
@(posedge clk);
#1;data_in = testData6[596];
@(posedge clk);
#1;data_in = testData6[597];
@(posedge clk);
#1;data_in = testData6[598];
@(posedge clk);
#1;data_in = testData6[599];
@(posedge clk);
#1;data_in = testData6[600];
@(posedge clk);
#1;data_in = testData6[601];
@(posedge clk);
#1;data_in = testData6[602];
@(posedge clk);
#1;data_in = testData6[603];
@(posedge clk);
#1;data_in = testData6[604];
@(posedge clk);
#1;data_in = testData6[605];
@(posedge clk);
#1;data_in = testData6[606];
@(posedge clk);
#1;data_in = testData6[607];
@(posedge clk);
#1;data_in = testData6[608];
@(posedge clk);
#1;data_in = testData6[609];
@(posedge clk);
#1;data_in = testData6[610];
@(posedge clk);
#1;data_in = testData6[611];
@(posedge clk);
#1;data_in = testData6[612];
@(posedge clk);
#1;data_in = testData6[613];
@(posedge clk);
#1;data_in = testData6[614];
@(posedge clk);
#1;data_in = testData6[615];
@(posedge clk);
#1;data_in = testData6[616];
@(posedge clk);
#1;data_in = testData6[617];
@(posedge clk);
#1;data_in = testData6[618];
@(posedge clk);
#1;data_in = testData6[619];
@(posedge clk);
#1;data_in = testData6[620];
@(posedge clk);
#1;data_in = testData6[621];
@(posedge clk);
#1;data_in = testData6[622];
@(posedge clk);
#1;data_in = testData6[623];
@(posedge clk);
#1;data_in = testData6[624];
@(posedge clk);
#1;data_in = testData6[625];
@(posedge clk);
#1;data_in = testData6[626];
@(posedge clk);
#1;data_in = testData6[627];
@(posedge clk);
#1;data_in = testData6[628];
@(posedge clk);
#1;data_in = testData6[629];
@(posedge clk);
#1;data_in = testData6[630];
@(posedge clk);
#1;data_in = testData6[631];
@(posedge clk);
#1;data_in = testData6[632];
@(posedge clk);
#1;data_in = testData6[633];
@(posedge clk);
#1;data_in = testData6[634];
@(posedge clk);
#1;data_in = testData6[635];
@(posedge clk);
#1;data_in = testData6[636];
@(posedge clk);
#1;data_in = testData6[637];
@(posedge clk);
#1;data_in = testData6[638];
@(posedge clk);
#1;data_in = testData6[639];
@(posedge clk);
#1;data_in = testData6[640];
@(posedge clk);
#1;data_in = testData6[641];
@(posedge clk);
#1;data_in = testData6[642];
@(posedge clk);
#1;data_in = testData6[643];
@(posedge clk);
#1;data_in = testData6[644];
@(posedge clk);
#1;data_in = testData6[645];
@(posedge clk);
#1;data_in = testData6[646];
@(posedge clk);
#1;data_in = testData6[647];
@(posedge clk);
#1;data_in = testData6[648];
@(posedge clk);
#1;data_in = testData6[649];
@(posedge clk);
#1;data_in = testData6[650];
@(posedge clk);
#1;data_in = testData6[651];
@(posedge clk);
#1;data_in = testData6[652];
@(posedge clk);
#1;data_in = testData6[653];
@(posedge clk);
#1;data_in = testData6[654];
@(posedge clk);
#1;data_in = testData6[655];
@(posedge clk);
#1;data_in = testData6[656];
@(posedge clk);
#1;data_in = testData6[657];
@(posedge clk);
#1;data_in = testData6[658];
@(posedge clk);
#1;data_in = testData6[659];
@(posedge clk);
#1;data_in = testData6[660];
@(posedge clk);
#1;data_in = testData6[661];
@(posedge clk);
#1;data_in = testData6[662];
@(posedge clk);
#1;data_in = testData6[663];
@(posedge clk);
#1;data_in = testData6[664];
@(posedge clk);
#1;data_in = testData6[665];
@(posedge clk);
#1;data_in = testData6[666];
@(posedge clk);
#1;data_in = testData6[667];
@(posedge clk);
#1;data_in = testData6[668];
@(posedge clk);
#1;data_in = testData6[669];
@(posedge clk);
#1;data_in = testData6[670];
@(posedge clk);
#1;data_in = testData6[671];
@(posedge clk);
#1;data_in = testData6[672];
@(posedge clk);
#1;data_in = testData6[673];
@(posedge clk);
#1;data_in = testData6[674];
@(posedge clk);
#1;data_in = testData6[675];
@(posedge clk);
#1;data_in = testData6[676];
@(posedge clk);
#1;data_in = testData6[677];
@(posedge clk);
#1;data_in = testData6[678];
@(posedge clk);
#1;data_in = testData6[679];
@(posedge clk);
#1;data_in = testData6[680];
@(posedge clk);
#1;data_in = testData6[681];
@(posedge clk);
#1;data_in = testData6[682];
@(posedge clk);
#1;data_in = testData6[683];
@(posedge clk);
#1;data_in = testData6[684];
@(posedge clk);
#1;data_in = testData6[685];
@(posedge clk);
#1;data_in = testData6[686];
@(posedge clk);
#1;data_in = testData6[687];
@(posedge clk);
#1;data_in = testData6[688];
@(posedge clk);
#1;data_in = testData6[689];
@(posedge clk);
#1;data_in = testData6[690];
@(posedge clk);
#1;data_in = testData6[691];
@(posedge clk);
#1;data_in = testData6[692];
@(posedge clk);
#1;data_in = testData6[693];
@(posedge clk);
#1;data_in = testData6[694];
@(posedge clk);
#1;data_in = testData6[695];
@(posedge clk);
#1;data_in = testData6[696];
@(posedge clk);
#1;data_in = testData6[697];
@(posedge clk);
#1;data_in = testData6[698];
@(posedge clk);
#1;data_in = testData6[699];
@(posedge clk);
#1;data_in = testData6[700];
@(posedge clk);
#1;data_in = testData6[701];
@(posedge clk);
#1;data_in = testData6[702];
@(posedge clk);
#1;data_in = testData6[703];
@(posedge clk);
#1;data_in = testData6[704];
@(posedge clk);
#1;data_in = testData6[705];
@(posedge clk);
#1;data_in = testData6[706];
@(posedge clk);
#1;data_in = testData6[707];
@(posedge clk);
#1;data_in = testData6[708];
@(posedge clk);
#1;data_in = testData6[709];
@(posedge clk);
#1;data_in = testData6[710];
@(posedge clk);
#1;data_in = testData6[711];
@(posedge clk);
#1;data_in = testData6[712];
@(posedge clk);
#1;data_in = testData6[713];
@(posedge clk);
#1;data_in = testData6[714];
@(posedge clk);
#1;data_in = testData6[715];
@(posedge clk);
#1;data_in = testData6[716];
@(posedge clk);
#1;data_in = testData6[717];
@(posedge clk);
#1;data_in = testData6[718];
@(posedge clk);
#1;data_in = testData6[719];
@(posedge clk);
#1;data_in = testData6[720];
@(posedge clk);
#1;data_in = testData6[721];
@(posedge clk);
#1;data_in = testData6[722];
@(posedge clk);
#1;data_in = testData6[723];
@(posedge clk);
#1;data_in = testData6[724];
@(posedge clk);
#1;data_in = testData6[725];
@(posedge clk);
#1;data_in = testData6[726];
@(posedge clk);
#1;data_in = testData6[727];
@(posedge clk);
#1;data_in = testData6[728];
@(posedge clk);
#1;data_in = testData6[729];
@(posedge clk);
#1;data_in = testData6[730];
@(posedge clk);
#1;data_in = testData6[731];
@(posedge clk);
#1;data_in = testData6[732];
@(posedge clk);
#1;data_in = testData6[733];
@(posedge clk);
#1;data_in = testData6[734];
@(posedge clk);
#1;data_in = testData6[735];
@(posedge clk);
#1;data_in = testData6[736];
@(posedge clk);
#1;data_in = testData6[737];
@(posedge clk);
#1;data_in = testData6[738];
@(posedge clk);
#1;data_in = testData6[739];
@(posedge clk);
#1;data_in = testData6[740];
@(posedge clk);
#1;data_in = testData6[741];
@(posedge clk);
#1;data_in = testData6[742];
@(posedge clk);
#1;data_in = testData6[743];
@(posedge clk);
#1;data_in = testData6[744];
@(posedge clk);
#1;data_in = testData6[745];
@(posedge clk);
#1;data_in = testData6[746];
@(posedge clk);
#1;data_in = testData6[747];
@(posedge clk);
#1;data_in = testData6[748];
@(posedge clk);
#1;data_in = testData6[749];
@(posedge clk);
#1;data_in = testData6[750];
@(posedge clk);
#1;data_in = testData6[751];
@(posedge clk);
#1;data_in = testData6[752];
@(posedge clk);
#1;data_in = testData6[753];
@(posedge clk);
#1;data_in = testData6[754];
@(posedge clk);
#1;data_in = testData6[755];
@(posedge clk);
#1;data_in = testData6[756];
@(posedge clk);
#1;data_in = testData6[757];
@(posedge clk);
#1;data_in = testData6[758];
@(posedge clk);
#1;data_in = testData6[759];
@(posedge clk);
#1;data_in = testData6[760];
@(posedge clk);
#1;data_in = testData6[761];
@(posedge clk);
#1;data_in = testData6[762];
@(posedge clk);
#1;data_in = testData6[763];
@(posedge clk);
#1;data_in = testData6[764];
@(posedge clk);
#1;data_in = testData6[765];
@(posedge clk);
#1;data_in = testData6[766];
@(posedge clk);
#1;data_in = testData6[767];
@(posedge clk);
#1;data_in = testData6[768];
@(posedge clk);
#1;data_in = testData6[769];
@(posedge clk);
#1;data_in = testData6[770];
@(posedge clk);
#1;data_in = testData6[771];
@(posedge clk);
#1;data_in = testData6[772];
@(posedge clk);
#1;data_in = testData6[773];
@(posedge clk);
#1;data_in = testData6[774];
@(posedge clk);
#1;data_in = testData6[775];
@(posedge clk);
#1;data_in = testData6[776];
@(posedge clk);
#1;data_in = testData6[777];
@(posedge clk);
#1;data_in = testData6[778];
@(posedge clk);
#1;data_in = testData6[779];
@(posedge clk);
#1;data_in = testData6[780];
@(posedge clk);
#1;data_in = testData6[781];
@(posedge clk);
#1;data_in = testData6[782];
@(posedge clk);
#1;data_in = testData6[783];
@(posedge clk);
#1;data_in = testData6[784];
@(posedge clk);
#1;data_in = testData6[785];
@(posedge clk);
#1;data_in = testData6[786];
@(posedge clk);
#1;data_in = testData6[787];
@(posedge clk);
#1;data_in = testData6[788];
@(posedge clk);
#1;data_in = testData6[789];
@(posedge clk);
#1;data_in = testData6[790];
@(posedge clk);
#1;data_in = testData6[791];
@(posedge clk);
#1;data_in = testData6[792];
@(posedge clk);
#1;data_in = testData6[793];
@(posedge clk);
#1;data_in = testData6[794];
@(posedge clk);
#1;data_in = testData6[795];
@(posedge clk);
#1;data_in = testData6[796];
@(posedge clk);
#1;data_in = testData6[797];
@(posedge clk);
#1;data_in = testData6[798];
@(posedge clk);
#1;data_in = testData6[799];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[800]; 
@(posedge clk);
#1;data_in = testData6[801];
@(posedge clk);
#1;data_in = testData6[802];
@(posedge clk);
#1;data_in = testData6[803];
@(posedge clk);
#1;data_in = testData6[804];
@(posedge clk);
#1;data_in = testData6[805];
@(posedge clk);
#1;data_in = testData6[806];
@(posedge clk);
#1;data_in = testData6[807];
@(posedge clk);
#1;data_in = testData6[808];
@(posedge clk);
#1;data_in = testData6[809];
@(posedge clk);
#1;data_in = testData6[810];
@(posedge clk);
#1;data_in = testData6[811];
@(posedge clk);
#1;data_in = testData6[812];
@(posedge clk);
#1;data_in = testData6[813];
@(posedge clk);
#1;data_in = testData6[814];
@(posedge clk);
#1;data_in = testData6[815];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[816];
@(posedge clk);
#1;data_in = testData6[817];
@(posedge clk);
#1;data_in = testData6[818];
@(posedge clk);
#1;data_in = testData6[819];
@(posedge clk);
#1;data_in = testData6[820];
@(posedge clk);
#1;data_in = testData6[821];
@(posedge clk);
#1;data_in = testData6[822];
@(posedge clk);
#1;data_in = testData6[823];
@(posedge clk);
#1;data_in = testData6[824];
@(posedge clk);
#1;data_in = testData6[825];
@(posedge clk);
#1;data_in = testData6[826];
@(posedge clk);
#1;data_in = testData6[827];
@(posedge clk);
#1;data_in = testData6[828];
@(posedge clk);
#1;data_in = testData6[829];
@(posedge clk);
#1;data_in = testData6[830];
@(posedge clk);
#1;data_in = testData6[831];
@(posedge clk);
#1;data_in = testData6[832];
@(posedge clk);
#1;data_in = testData6[833];
@(posedge clk);
#1;data_in = testData6[834];
@(posedge clk);
#1;data_in = testData6[835];
@(posedge clk);
#1;data_in = testData6[836];
@(posedge clk);
#1;data_in = testData6[837];
@(posedge clk);
#1;data_in = testData6[838];
@(posedge clk);
#1;data_in = testData6[839];
@(posedge clk);
#1;data_in = testData6[840];
@(posedge clk);
#1;data_in = testData6[841];
@(posedge clk);
#1;data_in = testData6[842];
@(posedge clk);
#1;data_in = testData6[843];
@(posedge clk);
#1;data_in = testData6[844];
@(posedge clk);
#1;data_in = testData6[845];
@(posedge clk);
#1;data_in = testData6[846];
@(posedge clk);
#1;data_in = testData6[847];
@(posedge clk);
#1;data_in = testData6[848];
@(posedge clk);
#1;data_in = testData6[849];
@(posedge clk);
#1;data_in = testData6[850];
@(posedge clk);
#1;data_in = testData6[851];
@(posedge clk);
#1;data_in = testData6[852];
@(posedge clk);
#1;data_in = testData6[853];
@(posedge clk);
#1;data_in = testData6[854];
@(posedge clk);
#1;data_in = testData6[855];
@(posedge clk);
#1;data_in = testData6[856];
@(posedge clk);
#1;data_in = testData6[857];
@(posedge clk);
#1;data_in = testData6[858];
@(posedge clk);
#1;data_in = testData6[859];
@(posedge clk);
#1;data_in = testData6[860];
@(posedge clk);
#1;data_in = testData6[861];
@(posedge clk);
#1;data_in = testData6[862];
@(posedge clk);
#1;data_in = testData6[863];
@(posedge clk);
#1;data_in = testData6[864];
@(posedge clk);
#1;data_in = testData6[865];
@(posedge clk);
#1;data_in = testData6[866];
@(posedge clk);
#1;data_in = testData6[867];
@(posedge clk);
#1;data_in = testData6[868];
@(posedge clk);
#1;data_in = testData6[869];
@(posedge clk);
#1;data_in = testData6[870];
@(posedge clk);
#1;data_in = testData6[871];
@(posedge clk);
#1;data_in = testData6[872];
@(posedge clk);
#1;data_in = testData6[873];
@(posedge clk);
#1;data_in = testData6[874];
@(posedge clk);
#1;data_in = testData6[875];
@(posedge clk);
#1;data_in = testData6[876];
@(posedge clk);
#1;data_in = testData6[877];
@(posedge clk);
#1;data_in = testData6[878];
@(posedge clk);
#1;data_in = testData6[879];
@(posedge clk);
#1;data_in = testData6[880];
@(posedge clk);
#1;data_in = testData6[881];
@(posedge clk);
#1;data_in = testData6[882];
@(posedge clk);
#1;data_in = testData6[883];
@(posedge clk);
#1;data_in = testData6[884];
@(posedge clk);
#1;data_in = testData6[885];
@(posedge clk);
#1;data_in = testData6[886];
@(posedge clk);
#1;data_in = testData6[887];
@(posedge clk);
#1;data_in = testData6[888];
@(posedge clk);
#1;data_in = testData6[889];
@(posedge clk);
#1;data_in = testData6[890];
@(posedge clk);
#1;data_in = testData6[891];
@(posedge clk);
#1;data_in = testData6[892];
@(posedge clk);
#1;data_in = testData6[893];
@(posedge clk);
#1;data_in = testData6[894];
@(posedge clk);
#1;data_in = testData6[895];
@(posedge clk);
#1;data_in = testData6[896];
@(posedge clk);
#1;data_in = testData6[897];
@(posedge clk);
#1;data_in = testData6[898];
@(posedge clk);
#1;data_in = testData6[899];
@(posedge clk);
#1;data_in = testData6[900];
@(posedge clk);
#1;data_in = testData6[901];
@(posedge clk);
#1;data_in = testData6[902];
@(posedge clk);
#1;data_in = testData6[903];
@(posedge clk);
#1;data_in = testData6[904];
@(posedge clk);
#1;data_in = testData6[905];
@(posedge clk);
#1;data_in = testData6[906];
@(posedge clk);
#1;data_in = testData6[907];
@(posedge clk);
#1;data_in = testData6[908];
@(posedge clk);
#1;data_in = testData6[909];
@(posedge clk);
#1;data_in = testData6[910];
@(posedge clk);
#1;data_in = testData6[911];
@(posedge clk);
#1;data_in = testData6[912];
@(posedge clk);
#1;data_in = testData6[913];
@(posedge clk);
#1;data_in = testData6[914];
@(posedge clk);
#1;data_in = testData6[915];
@(posedge clk);
#1;data_in = testData6[916];
@(posedge clk);
#1;data_in = testData6[917];
@(posedge clk);
#1;data_in = testData6[918];
@(posedge clk);
#1;data_in = testData6[919];
@(posedge clk);
#1;data_in = testData6[920];
@(posedge clk);
#1;data_in = testData6[921];
@(posedge clk);
#1;data_in = testData6[922];
@(posedge clk);
#1;data_in = testData6[923];
@(posedge clk);
#1;data_in = testData6[924];
@(posedge clk);
#1;data_in = testData6[925];
@(posedge clk);
#1;data_in = testData6[926];
@(posedge clk);
#1;data_in = testData6[927];
@(posedge clk);
#1;data_in = testData6[928];
@(posedge clk);
#1;data_in = testData6[929];
@(posedge clk);
#1;data_in = testData6[930];
@(posedge clk);
#1;data_in = testData6[931];
@(posedge clk);
#1;data_in = testData6[932];
@(posedge clk);
#1;data_in = testData6[933];
@(posedge clk);
#1;data_in = testData6[934];
@(posedge clk);
#1;data_in = testData6[935];
@(posedge clk);
#1;data_in = testData6[936];
@(posedge clk);
#1;data_in = testData6[937];
@(posedge clk);
#1;data_in = testData6[938];
@(posedge clk);
#1;data_in = testData6[939];
@(posedge clk);
#1;data_in = testData6[940];
@(posedge clk);
#1;data_in = testData6[941];
@(posedge clk);
#1;data_in = testData6[942];
@(posedge clk);
#1;data_in = testData6[943];
@(posedge clk);
#1;data_in = testData6[944];
@(posedge clk);
#1;data_in = testData6[945];
@(posedge clk);
#1;data_in = testData6[946];
@(posedge clk);
#1;data_in = testData6[947];
@(posedge clk);
#1;data_in = testData6[948];
@(posedge clk);
#1;data_in = testData6[949];
@(posedge clk);
#1;data_in = testData6[950];
@(posedge clk);
#1;data_in = testData6[951];
@(posedge clk);
#1;data_in = testData6[952];
@(posedge clk);
#1;data_in = testData6[953];
@(posedge clk);
#1;data_in = testData6[954];
@(posedge clk);
#1;data_in = testData6[955];
@(posedge clk);
#1;data_in = testData6[956];
@(posedge clk);
#1;data_in = testData6[957];
@(posedge clk);
#1;data_in = testData6[958];
@(posedge clk);
#1;data_in = testData6[959];
@(posedge clk);
#1;data_in = testData6[960];
@(posedge clk);
#1;data_in = testData6[961];
@(posedge clk);
#1;data_in = testData6[962];
@(posedge clk);
#1;data_in = testData6[963];
@(posedge clk);
#1;data_in = testData6[964];
@(posedge clk);
#1;data_in = testData6[965];
@(posedge clk);
#1;data_in = testData6[966];
@(posedge clk);
#1;data_in = testData6[967];
@(posedge clk);
#1;data_in = testData6[968];
@(posedge clk);
#1;data_in = testData6[969];
@(posedge clk);
#1;data_in = testData6[970];
@(posedge clk);
#1;data_in = testData6[971];
@(posedge clk);
#1;data_in = testData6[972];
@(posedge clk);
#1;data_in = testData6[973];
@(posedge clk);
#1;data_in = testData6[974];
@(posedge clk);
#1;data_in = testData6[975];
@(posedge clk);
#1;data_in = testData6[976];
@(posedge clk);
#1;data_in = testData6[977];
@(posedge clk);
#1;data_in = testData6[978];
@(posedge clk);
#1;data_in = testData6[979];
@(posedge clk);
#1;data_in = testData6[980];
@(posedge clk);
#1;data_in = testData6[981];
@(posedge clk);
#1;data_in = testData6[982];
@(posedge clk);
#1;data_in = testData6[983];
@(posedge clk);
#1;data_in = testData6[984];
@(posedge clk);
#1;data_in = testData6[985];
@(posedge clk);
#1;data_in = testData6[986];
@(posedge clk);
#1;data_in = testData6[987];
@(posedge clk);
#1;data_in = testData6[988];
@(posedge clk);
#1;data_in = testData6[989];
@(posedge clk);
#1;data_in = testData6[990];
@(posedge clk);
#1;data_in = testData6[991];
@(posedge clk);
#1;data_in = testData6[992];
@(posedge clk);
#1;data_in = testData6[993];
@(posedge clk);
#1;data_in = testData6[994];
@(posedge clk);
#1;data_in = testData6[995];
@(posedge clk);
#1;data_in = testData6[996];
@(posedge clk);
#1;data_in = testData6[997];
@(posedge clk);
#1;data_in = testData6[998];
@(posedge clk);
#1;data_in = testData6[999];
@(posedge clk);
#1;data_in = testData6[1000];
@(posedge clk);
#1;data_in = testData6[1001];
@(posedge clk);
#1;data_in = testData6[1002];
@(posedge clk);
#1;data_in = testData6[1003];
@(posedge clk);
#1;data_in = testData6[1004];
@(posedge clk);
#1;data_in = testData6[1005];
@(posedge clk);
#1;data_in = testData6[1006];
@(posedge clk);
#1;data_in = testData6[1007];
@(posedge clk);
#1;data_in = testData6[1008];
@(posedge clk);
#1;data_in = testData6[1009];
@(posedge clk);
#1;data_in = testData6[1010];
@(posedge clk);
#1;data_in = testData6[1011];
@(posedge clk);
#1;data_in = testData6[1012];
@(posedge clk);
#1;data_in = testData6[1013];
@(posedge clk);
#1;data_in = testData6[1014];
@(posedge clk);
#1;data_in = testData6[1015];
@(posedge clk);
#1;data_in = testData6[1016];
@(posedge clk);
#1;data_in = testData6[1017];
@(posedge clk);
#1;data_in = testData6[1018];
@(posedge clk);
#1;data_in = testData6[1019];
@(posedge clk);
#1;data_in = testData6[1020];
@(posedge clk);
#1;data_in = testData6[1021];
@(posedge clk);
#1;data_in = testData6[1022];
@(posedge clk);
#1;data_in = testData6[1023];
@(posedge clk);
#1;data_in = testData6[1024];
@(posedge clk);
#1;data_in = testData6[1025];
@(posedge clk);
#1;data_in = testData6[1026];
@(posedge clk);
#1;data_in = testData6[1027];
@(posedge clk);
#1;data_in = testData6[1028];
@(posedge clk);
#1;data_in = testData6[1029];
@(posedge clk);
#1;data_in = testData6[1030];
@(posedge clk);
#1;data_in = testData6[1031];
@(posedge clk);
#1;data_in = testData6[1032];
@(posedge clk);
#1;data_in = testData6[1033];
@(posedge clk);
#1;data_in = testData6[1034];
@(posedge clk);
#1;data_in = testData6[1035];
@(posedge clk);
#1;data_in = testData6[1036];
@(posedge clk);
#1;data_in = testData6[1037];
@(posedge clk);
#1;data_in = testData6[1038];
@(posedge clk);
#1;data_in = testData6[1039];
@(posedge clk);
#1;data_in = testData6[1040];
@(posedge clk);
#1;data_in = testData6[1041];
@(posedge clk);
#1;data_in = testData6[1042];
@(posedge clk);
#1;data_in = testData6[1043];
@(posedge clk);
#1;data_in = testData6[1044];
@(posedge clk);
#1;data_in = testData6[1045];
@(posedge clk);
#1;data_in = testData6[1046];
@(posedge clk);
#1;data_in = testData6[1047];
@(posedge clk);
#1;data_in = testData6[1048];
@(posedge clk);
#1;data_in = testData6[1049];
@(posedge clk);
#1;data_in = testData6[1050];
@(posedge clk);
#1;data_in = testData6[1051];
@(posedge clk);
#1;data_in = testData6[1052];
@(posedge clk);
#1;data_in = testData6[1053];
@(posedge clk);
#1;data_in = testData6[1054];
@(posedge clk);
#1;data_in = testData6[1055];
@(posedge clk);
#1;data_in = testData6[1056];
@(posedge clk);
#1;data_in = testData6[1057];
@(posedge clk);
#1;data_in = testData6[1058];
@(posedge clk);
#1;data_in = testData6[1059];
@(posedge clk);
#1;data_in = testData6[1060];
@(posedge clk);
#1;data_in = testData6[1061];
@(posedge clk);
#1;data_in = testData6[1062];
@(posedge clk);
#1;data_in = testData6[1063];
@(posedge clk);
#1;data_in = testData6[1064];
@(posedge clk);
#1;data_in = testData6[1065];
@(posedge clk);
#1;data_in = testData6[1066];
@(posedge clk);
#1;data_in = testData6[1067];
@(posedge clk);
#1;data_in = testData6[1068];
@(posedge clk);
#1;data_in = testData6[1069];
@(posedge clk);
#1;data_in = testData6[1070];
@(posedge clk);
#1;data_in = testData6[1071];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1072]; 
@(posedge clk);
#1;data_in = testData6[1073];
@(posedge clk);
#1;data_in = testData6[1074];
@(posedge clk);
#1;data_in = testData6[1075];
@(posedge clk);
#1;data_in = testData6[1076];
@(posedge clk);
#1;data_in = testData6[1077];
@(posedge clk);
#1;data_in = testData6[1078];
@(posedge clk);
#1;data_in = testData6[1079];
@(posedge clk);
#1;data_in = testData6[1080];
@(posedge clk);
#1;data_in = testData6[1081];
@(posedge clk);
#1;data_in = testData6[1082];
@(posedge clk);
#1;data_in = testData6[1083];
@(posedge clk);
#1;data_in = testData6[1084];
@(posedge clk);
#1;data_in = testData6[1085];
@(posedge clk);
#1;data_in = testData6[1086];
@(posedge clk);
#1;data_in = testData6[1087];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1088];
@(posedge clk);
#1;data_in = testData6[1089];
@(posedge clk);
#1;data_in = testData6[1090];
@(posedge clk);
#1;data_in = testData6[1091];
@(posedge clk);
#1;data_in = testData6[1092];
@(posedge clk);
#1;data_in = testData6[1093];
@(posedge clk);
#1;data_in = testData6[1094];
@(posedge clk);
#1;data_in = testData6[1095];
@(posedge clk);
#1;data_in = testData6[1096];
@(posedge clk);
#1;data_in = testData6[1097];
@(posedge clk);
#1;data_in = testData6[1098];
@(posedge clk);
#1;data_in = testData6[1099];
@(posedge clk);
#1;data_in = testData6[1100];
@(posedge clk);
#1;data_in = testData6[1101];
@(posedge clk);
#1;data_in = testData6[1102];
@(posedge clk);
#1;data_in = testData6[1103];
@(posedge clk);
#1;data_in = testData6[1104];
@(posedge clk);
#1;data_in = testData6[1105];
@(posedge clk);
#1;data_in = testData6[1106];
@(posedge clk);
#1;data_in = testData6[1107];
@(posedge clk);
#1;data_in = testData6[1108];
@(posedge clk);
#1;data_in = testData6[1109];
@(posedge clk);
#1;data_in = testData6[1110];
@(posedge clk);
#1;data_in = testData6[1111];
@(posedge clk);
#1;data_in = testData6[1112];
@(posedge clk);
#1;data_in = testData6[1113];
@(posedge clk);
#1;data_in = testData6[1114];
@(posedge clk);
#1;data_in = testData6[1115];
@(posedge clk);
#1;data_in = testData6[1116];
@(posedge clk);
#1;data_in = testData6[1117];
@(posedge clk);
#1;data_in = testData6[1118];
@(posedge clk);
#1;data_in = testData6[1119];
@(posedge clk);
#1;data_in = testData6[1120];
@(posedge clk);
#1;data_in = testData6[1121];
@(posedge clk);
#1;data_in = testData6[1122];
@(posedge clk);
#1;data_in = testData6[1123];
@(posedge clk);
#1;data_in = testData6[1124];
@(posedge clk);
#1;data_in = testData6[1125];
@(posedge clk);
#1;data_in = testData6[1126];
@(posedge clk);
#1;data_in = testData6[1127];
@(posedge clk);
#1;data_in = testData6[1128];
@(posedge clk);
#1;data_in = testData6[1129];
@(posedge clk);
#1;data_in = testData6[1130];
@(posedge clk);
#1;data_in = testData6[1131];
@(posedge clk);
#1;data_in = testData6[1132];
@(posedge clk);
#1;data_in = testData6[1133];
@(posedge clk);
#1;data_in = testData6[1134];
@(posedge clk);
#1;data_in = testData6[1135];
@(posedge clk);
#1;data_in = testData6[1136];
@(posedge clk);
#1;data_in = testData6[1137];
@(posedge clk);
#1;data_in = testData6[1138];
@(posedge clk);
#1;data_in = testData6[1139];
@(posedge clk);
#1;data_in = testData6[1140];
@(posedge clk);
#1;data_in = testData6[1141];
@(posedge clk);
#1;data_in = testData6[1142];
@(posedge clk);
#1;data_in = testData6[1143];
@(posedge clk);
#1;data_in = testData6[1144];
@(posedge clk);
#1;data_in = testData6[1145];
@(posedge clk);
#1;data_in = testData6[1146];
@(posedge clk);
#1;data_in = testData6[1147];
@(posedge clk);
#1;data_in = testData6[1148];
@(posedge clk);
#1;data_in = testData6[1149];
@(posedge clk);
#1;data_in = testData6[1150];
@(posedge clk);
#1;data_in = testData6[1151];
@(posedge clk);
#1;data_in = testData6[1152];
@(posedge clk);
#1;data_in = testData6[1153];
@(posedge clk);
#1;data_in = testData6[1154];
@(posedge clk);
#1;data_in = testData6[1155];
@(posedge clk);
#1;data_in = testData6[1156];
@(posedge clk);
#1;data_in = testData6[1157];
@(posedge clk);
#1;data_in = testData6[1158];
@(posedge clk);
#1;data_in = testData6[1159];
@(posedge clk);
#1;data_in = testData6[1160];
@(posedge clk);
#1;data_in = testData6[1161];
@(posedge clk);
#1;data_in = testData6[1162];
@(posedge clk);
#1;data_in = testData6[1163];
@(posedge clk);
#1;data_in = testData6[1164];
@(posedge clk);
#1;data_in = testData6[1165];
@(posedge clk);
#1;data_in = testData6[1166];
@(posedge clk);
#1;data_in = testData6[1167];
@(posedge clk);
#1;data_in = testData6[1168];
@(posedge clk);
#1;data_in = testData6[1169];
@(posedge clk);
#1;data_in = testData6[1170];
@(posedge clk);
#1;data_in = testData6[1171];
@(posedge clk);
#1;data_in = testData6[1172];
@(posedge clk);
#1;data_in = testData6[1173];
@(posedge clk);
#1;data_in = testData6[1174];
@(posedge clk);
#1;data_in = testData6[1175];
@(posedge clk);
#1;data_in = testData6[1176];
@(posedge clk);
#1;data_in = testData6[1177];
@(posedge clk);
#1;data_in = testData6[1178];
@(posedge clk);
#1;data_in = testData6[1179];
@(posedge clk);
#1;data_in = testData6[1180];
@(posedge clk);
#1;data_in = testData6[1181];
@(posedge clk);
#1;data_in = testData6[1182];
@(posedge clk);
#1;data_in = testData6[1183];
@(posedge clk);
#1;data_in = testData6[1184];
@(posedge clk);
#1;data_in = testData6[1185];
@(posedge clk);
#1;data_in = testData6[1186];
@(posedge clk);
#1;data_in = testData6[1187];
@(posedge clk);
#1;data_in = testData6[1188];
@(posedge clk);
#1;data_in = testData6[1189];
@(posedge clk);
#1;data_in = testData6[1190];
@(posedge clk);
#1;data_in = testData6[1191];
@(posedge clk);
#1;data_in = testData6[1192];
@(posedge clk);
#1;data_in = testData6[1193];
@(posedge clk);
#1;data_in = testData6[1194];
@(posedge clk);
#1;data_in = testData6[1195];
@(posedge clk);
#1;data_in = testData6[1196];
@(posedge clk);
#1;data_in = testData6[1197];
@(posedge clk);
#1;data_in = testData6[1198];
@(posedge clk);
#1;data_in = testData6[1199];
@(posedge clk);
#1;data_in = testData6[1200];
@(posedge clk);
#1;data_in = testData6[1201];
@(posedge clk);
#1;data_in = testData6[1202];
@(posedge clk);
#1;data_in = testData6[1203];
@(posedge clk);
#1;data_in = testData6[1204];
@(posedge clk);
#1;data_in = testData6[1205];
@(posedge clk);
#1;data_in = testData6[1206];
@(posedge clk);
#1;data_in = testData6[1207];
@(posedge clk);
#1;data_in = testData6[1208];
@(posedge clk);
#1;data_in = testData6[1209];
@(posedge clk);
#1;data_in = testData6[1210];
@(posedge clk);
#1;data_in = testData6[1211];
@(posedge clk);
#1;data_in = testData6[1212];
@(posedge clk);
#1;data_in = testData6[1213];
@(posedge clk);
#1;data_in = testData6[1214];
@(posedge clk);
#1;data_in = testData6[1215];
@(posedge clk);
#1;data_in = testData6[1216];
@(posedge clk);
#1;data_in = testData6[1217];
@(posedge clk);
#1;data_in = testData6[1218];
@(posedge clk);
#1;data_in = testData6[1219];
@(posedge clk);
#1;data_in = testData6[1220];
@(posedge clk);
#1;data_in = testData6[1221];
@(posedge clk);
#1;data_in = testData6[1222];
@(posedge clk);
#1;data_in = testData6[1223];
@(posedge clk);
#1;data_in = testData6[1224];
@(posedge clk);
#1;data_in = testData6[1225];
@(posedge clk);
#1;data_in = testData6[1226];
@(posedge clk);
#1;data_in = testData6[1227];
@(posedge clk);
#1;data_in = testData6[1228];
@(posedge clk);
#1;data_in = testData6[1229];
@(posedge clk);
#1;data_in = testData6[1230];
@(posedge clk);
#1;data_in = testData6[1231];
@(posedge clk);
#1;data_in = testData6[1232];
@(posedge clk);
#1;data_in = testData6[1233];
@(posedge clk);
#1;data_in = testData6[1234];
@(posedge clk);
#1;data_in = testData6[1235];
@(posedge clk);
#1;data_in = testData6[1236];
@(posedge clk);
#1;data_in = testData6[1237];
@(posedge clk);
#1;data_in = testData6[1238];
@(posedge clk);
#1;data_in = testData6[1239];
@(posedge clk);
#1;data_in = testData6[1240];
@(posedge clk);
#1;data_in = testData6[1241];
@(posedge clk);
#1;data_in = testData6[1242];
@(posedge clk);
#1;data_in = testData6[1243];
@(posedge clk);
#1;data_in = testData6[1244];
@(posedge clk);
#1;data_in = testData6[1245];
@(posedge clk);
#1;data_in = testData6[1246];
@(posedge clk);
#1;data_in = testData6[1247];
@(posedge clk);
#1;data_in = testData6[1248];
@(posedge clk);
#1;data_in = testData6[1249];
@(posedge clk);
#1;data_in = testData6[1250];
@(posedge clk);
#1;data_in = testData6[1251];
@(posedge clk);
#1;data_in = testData6[1252];
@(posedge clk);
#1;data_in = testData6[1253];
@(posedge clk);
#1;data_in = testData6[1254];
@(posedge clk);
#1;data_in = testData6[1255];
@(posedge clk);
#1;data_in = testData6[1256];
@(posedge clk);
#1;data_in = testData6[1257];
@(posedge clk);
#1;data_in = testData6[1258];
@(posedge clk);
#1;data_in = testData6[1259];
@(posedge clk);
#1;data_in = testData6[1260];
@(posedge clk);
#1;data_in = testData6[1261];
@(posedge clk);
#1;data_in = testData6[1262];
@(posedge clk);
#1;data_in = testData6[1263];
@(posedge clk);
#1;data_in = testData6[1264];
@(posedge clk);
#1;data_in = testData6[1265];
@(posedge clk);
#1;data_in = testData6[1266];
@(posedge clk);
#1;data_in = testData6[1267];
@(posedge clk);
#1;data_in = testData6[1268];
@(posedge clk);
#1;data_in = testData6[1269];
@(posedge clk);
#1;data_in = testData6[1270];
@(posedge clk);
#1;data_in = testData6[1271];
@(posedge clk);
#1;data_in = testData6[1272];
@(posedge clk);
#1;data_in = testData6[1273];
@(posedge clk);
#1;data_in = testData6[1274];
@(posedge clk);
#1;data_in = testData6[1275];
@(posedge clk);
#1;data_in = testData6[1276];
@(posedge clk);
#1;data_in = testData6[1277];
@(posedge clk);
#1;data_in = testData6[1278];
@(posedge clk);
#1;data_in = testData6[1279];
@(posedge clk);
#1;data_in = testData6[1280];
@(posedge clk);
#1;data_in = testData6[1281];
@(posedge clk);
#1;data_in = testData6[1282];
@(posedge clk);
#1;data_in = testData6[1283];
@(posedge clk);
#1;data_in = testData6[1284];
@(posedge clk);
#1;data_in = testData6[1285];
@(posedge clk);
#1;data_in = testData6[1286];
@(posedge clk);
#1;data_in = testData6[1287];
@(posedge clk);
#1;data_in = testData6[1288];
@(posedge clk);
#1;data_in = testData6[1289];
@(posedge clk);
#1;data_in = testData6[1290];
@(posedge clk);
#1;data_in = testData6[1291];
@(posedge clk);
#1;data_in = testData6[1292];
@(posedge clk);
#1;data_in = testData6[1293];
@(posedge clk);
#1;data_in = testData6[1294];
@(posedge clk);
#1;data_in = testData6[1295];
@(posedge clk);
#1;data_in = testData6[1296];
@(posedge clk);
#1;data_in = testData6[1297];
@(posedge clk);
#1;data_in = testData6[1298];
@(posedge clk);
#1;data_in = testData6[1299];
@(posedge clk);
#1;data_in = testData6[1300];
@(posedge clk);
#1;data_in = testData6[1301];
@(posedge clk);
#1;data_in = testData6[1302];
@(posedge clk);
#1;data_in = testData6[1303];
@(posedge clk);
#1;data_in = testData6[1304];
@(posedge clk);
#1;data_in = testData6[1305];
@(posedge clk);
#1;data_in = testData6[1306];
@(posedge clk);
#1;data_in = testData6[1307];
@(posedge clk);
#1;data_in = testData6[1308];
@(posedge clk);
#1;data_in = testData6[1309];
@(posedge clk);
#1;data_in = testData6[1310];
@(posedge clk);
#1;data_in = testData6[1311];
@(posedge clk);
#1;data_in = testData6[1312];
@(posedge clk);
#1;data_in = testData6[1313];
@(posedge clk);
#1;data_in = testData6[1314];
@(posedge clk);
#1;data_in = testData6[1315];
@(posedge clk);
#1;data_in = testData6[1316];
@(posedge clk);
#1;data_in = testData6[1317];
@(posedge clk);
#1;data_in = testData6[1318];
@(posedge clk);
#1;data_in = testData6[1319];
@(posedge clk);
#1;data_in = testData6[1320];
@(posedge clk);
#1;data_in = testData6[1321];
@(posedge clk);
#1;data_in = testData6[1322];
@(posedge clk);
#1;data_in = testData6[1323];
@(posedge clk);
#1;data_in = testData6[1324];
@(posedge clk);
#1;data_in = testData6[1325];
@(posedge clk);
#1;data_in = testData6[1326];
@(posedge clk);
#1;data_in = testData6[1327];
@(posedge clk);
#1;data_in = testData6[1328];
@(posedge clk);
#1;data_in = testData6[1329];
@(posedge clk);
#1;data_in = testData6[1330];
@(posedge clk);
#1;data_in = testData6[1331];
@(posedge clk);
#1;data_in = testData6[1332];
@(posedge clk);
#1;data_in = testData6[1333];
@(posedge clk);
#1;data_in = testData6[1334];
@(posedge clk);
#1;data_in = testData6[1335];
@(posedge clk);
#1;data_in = testData6[1336];
@(posedge clk);
#1;data_in = testData6[1337];
@(posedge clk);
#1;data_in = testData6[1338];
@(posedge clk);
#1;data_in = testData6[1339];
@(posedge clk);
#1;data_in = testData6[1340];
@(posedge clk);
#1;data_in = testData6[1341];
@(posedge clk);
#1;data_in = testData6[1342];
@(posedge clk);
#1;data_in = testData6[1343];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1344]; 
@(posedge clk);
#1;data_in = testData6[1345];
@(posedge clk);
#1;data_in = testData6[1346];
@(posedge clk);
#1;data_in = testData6[1347];
@(posedge clk);
#1;data_in = testData6[1348];
@(posedge clk);
#1;data_in = testData6[1349];
@(posedge clk);
#1;data_in = testData6[1350];
@(posedge clk);
#1;data_in = testData6[1351];
@(posedge clk);
#1;data_in = testData6[1352];
@(posedge clk);
#1;data_in = testData6[1353];
@(posedge clk);
#1;data_in = testData6[1354];
@(posedge clk);
#1;data_in = testData6[1355];
@(posedge clk);
#1;data_in = testData6[1356];
@(posedge clk);
#1;data_in = testData6[1357];
@(posedge clk);
#1;data_in = testData6[1358];
@(posedge clk);
#1;data_in = testData6[1359];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1360];
@(posedge clk);
#1;data_in = testData6[1361];
@(posedge clk);
#1;data_in = testData6[1362];
@(posedge clk);
#1;data_in = testData6[1363];
@(posedge clk);
#1;data_in = testData6[1364];
@(posedge clk);
#1;data_in = testData6[1365];
@(posedge clk);
#1;data_in = testData6[1366];
@(posedge clk);
#1;data_in = testData6[1367];
@(posedge clk);
#1;data_in = testData6[1368];
@(posedge clk);
#1;data_in = testData6[1369];
@(posedge clk);
#1;data_in = testData6[1370];
@(posedge clk);
#1;data_in = testData6[1371];
@(posedge clk);
#1;data_in = testData6[1372];
@(posedge clk);
#1;data_in = testData6[1373];
@(posedge clk);
#1;data_in = testData6[1374];
@(posedge clk);
#1;data_in = testData6[1375];
@(posedge clk);
#1;data_in = testData6[1376];
@(posedge clk);
#1;data_in = testData6[1377];
@(posedge clk);
#1;data_in = testData6[1378];
@(posedge clk);
#1;data_in = testData6[1379];
@(posedge clk);
#1;data_in = testData6[1380];
@(posedge clk);
#1;data_in = testData6[1381];
@(posedge clk);
#1;data_in = testData6[1382];
@(posedge clk);
#1;data_in = testData6[1383];
@(posedge clk);
#1;data_in = testData6[1384];
@(posedge clk);
#1;data_in = testData6[1385];
@(posedge clk);
#1;data_in = testData6[1386];
@(posedge clk);
#1;data_in = testData6[1387];
@(posedge clk);
#1;data_in = testData6[1388];
@(posedge clk);
#1;data_in = testData6[1389];
@(posedge clk);
#1;data_in = testData6[1390];
@(posedge clk);
#1;data_in = testData6[1391];
@(posedge clk);
#1;data_in = testData6[1392];
@(posedge clk);
#1;data_in = testData6[1393];
@(posedge clk);
#1;data_in = testData6[1394];
@(posedge clk);
#1;data_in = testData6[1395];
@(posedge clk);
#1;data_in = testData6[1396];
@(posedge clk);
#1;data_in = testData6[1397];
@(posedge clk);
#1;data_in = testData6[1398];
@(posedge clk);
#1;data_in = testData6[1399];
@(posedge clk);
#1;data_in = testData6[1400];
@(posedge clk);
#1;data_in = testData6[1401];
@(posedge clk);
#1;data_in = testData6[1402];
@(posedge clk);
#1;data_in = testData6[1403];
@(posedge clk);
#1;data_in = testData6[1404];
@(posedge clk);
#1;data_in = testData6[1405];
@(posedge clk);
#1;data_in = testData6[1406];
@(posedge clk);
#1;data_in = testData6[1407];
@(posedge clk);
#1;data_in = testData6[1408];
@(posedge clk);
#1;data_in = testData6[1409];
@(posedge clk);
#1;data_in = testData6[1410];
@(posedge clk);
#1;data_in = testData6[1411];
@(posedge clk);
#1;data_in = testData6[1412];
@(posedge clk);
#1;data_in = testData6[1413];
@(posedge clk);
#1;data_in = testData6[1414];
@(posedge clk);
#1;data_in = testData6[1415];
@(posedge clk);
#1;data_in = testData6[1416];
@(posedge clk);
#1;data_in = testData6[1417];
@(posedge clk);
#1;data_in = testData6[1418];
@(posedge clk);
#1;data_in = testData6[1419];
@(posedge clk);
#1;data_in = testData6[1420];
@(posedge clk);
#1;data_in = testData6[1421];
@(posedge clk);
#1;data_in = testData6[1422];
@(posedge clk);
#1;data_in = testData6[1423];
@(posedge clk);
#1;data_in = testData6[1424];
@(posedge clk);
#1;data_in = testData6[1425];
@(posedge clk);
#1;data_in = testData6[1426];
@(posedge clk);
#1;data_in = testData6[1427];
@(posedge clk);
#1;data_in = testData6[1428];
@(posedge clk);
#1;data_in = testData6[1429];
@(posedge clk);
#1;data_in = testData6[1430];
@(posedge clk);
#1;data_in = testData6[1431];
@(posedge clk);
#1;data_in = testData6[1432];
@(posedge clk);
#1;data_in = testData6[1433];
@(posedge clk);
#1;data_in = testData6[1434];
@(posedge clk);
#1;data_in = testData6[1435];
@(posedge clk);
#1;data_in = testData6[1436];
@(posedge clk);
#1;data_in = testData6[1437];
@(posedge clk);
#1;data_in = testData6[1438];
@(posedge clk);
#1;data_in = testData6[1439];
@(posedge clk);
#1;data_in = testData6[1440];
@(posedge clk);
#1;data_in = testData6[1441];
@(posedge clk);
#1;data_in = testData6[1442];
@(posedge clk);
#1;data_in = testData6[1443];
@(posedge clk);
#1;data_in = testData6[1444];
@(posedge clk);
#1;data_in = testData6[1445];
@(posedge clk);
#1;data_in = testData6[1446];
@(posedge clk);
#1;data_in = testData6[1447];
@(posedge clk);
#1;data_in = testData6[1448];
@(posedge clk);
#1;data_in = testData6[1449];
@(posedge clk);
#1;data_in = testData6[1450];
@(posedge clk);
#1;data_in = testData6[1451];
@(posedge clk);
#1;data_in = testData6[1452];
@(posedge clk);
#1;data_in = testData6[1453];
@(posedge clk);
#1;data_in = testData6[1454];
@(posedge clk);
#1;data_in = testData6[1455];
@(posedge clk);
#1;data_in = testData6[1456];
@(posedge clk);
#1;data_in = testData6[1457];
@(posedge clk);
#1;data_in = testData6[1458];
@(posedge clk);
#1;data_in = testData6[1459];
@(posedge clk);
#1;data_in = testData6[1460];
@(posedge clk);
#1;data_in = testData6[1461];
@(posedge clk);
#1;data_in = testData6[1462];
@(posedge clk);
#1;data_in = testData6[1463];
@(posedge clk);
#1;data_in = testData6[1464];
@(posedge clk);
#1;data_in = testData6[1465];
@(posedge clk);
#1;data_in = testData6[1466];
@(posedge clk);
#1;data_in = testData6[1467];
@(posedge clk);
#1;data_in = testData6[1468];
@(posedge clk);
#1;data_in = testData6[1469];
@(posedge clk);
#1;data_in = testData6[1470];
@(posedge clk);
#1;data_in = testData6[1471];
@(posedge clk);
#1;data_in = testData6[1472];
@(posedge clk);
#1;data_in = testData6[1473];
@(posedge clk);
#1;data_in = testData6[1474];
@(posedge clk);
#1;data_in = testData6[1475];
@(posedge clk);
#1;data_in = testData6[1476];
@(posedge clk);
#1;data_in = testData6[1477];
@(posedge clk);
#1;data_in = testData6[1478];
@(posedge clk);
#1;data_in = testData6[1479];
@(posedge clk);
#1;data_in = testData6[1480];
@(posedge clk);
#1;data_in = testData6[1481];
@(posedge clk);
#1;data_in = testData6[1482];
@(posedge clk);
#1;data_in = testData6[1483];
@(posedge clk);
#1;data_in = testData6[1484];
@(posedge clk);
#1;data_in = testData6[1485];
@(posedge clk);
#1;data_in = testData6[1486];
@(posedge clk);
#1;data_in = testData6[1487];
@(posedge clk);
#1;data_in = testData6[1488];
@(posedge clk);
#1;data_in = testData6[1489];
@(posedge clk);
#1;data_in = testData6[1490];
@(posedge clk);
#1;data_in = testData6[1491];
@(posedge clk);
#1;data_in = testData6[1492];
@(posedge clk);
#1;data_in = testData6[1493];
@(posedge clk);
#1;data_in = testData6[1494];
@(posedge clk);
#1;data_in = testData6[1495];
@(posedge clk);
#1;data_in = testData6[1496];
@(posedge clk);
#1;data_in = testData6[1497];
@(posedge clk);
#1;data_in = testData6[1498];
@(posedge clk);
#1;data_in = testData6[1499];
@(posedge clk);
#1;data_in = testData6[1500];
@(posedge clk);
#1;data_in = testData6[1501];
@(posedge clk);
#1;data_in = testData6[1502];
@(posedge clk);
#1;data_in = testData6[1503];
@(posedge clk);
#1;data_in = testData6[1504];
@(posedge clk);
#1;data_in = testData6[1505];
@(posedge clk);
#1;data_in = testData6[1506];
@(posedge clk);
#1;data_in = testData6[1507];
@(posedge clk);
#1;data_in = testData6[1508];
@(posedge clk);
#1;data_in = testData6[1509];
@(posedge clk);
#1;data_in = testData6[1510];
@(posedge clk);
#1;data_in = testData6[1511];
@(posedge clk);
#1;data_in = testData6[1512];
@(posedge clk);
#1;data_in = testData6[1513];
@(posedge clk);
#1;data_in = testData6[1514];
@(posedge clk);
#1;data_in = testData6[1515];
@(posedge clk);
#1;data_in = testData6[1516];
@(posedge clk);
#1;data_in = testData6[1517];
@(posedge clk);
#1;data_in = testData6[1518];
@(posedge clk);
#1;data_in = testData6[1519];
@(posedge clk);
#1;data_in = testData6[1520];
@(posedge clk);
#1;data_in = testData6[1521];
@(posedge clk);
#1;data_in = testData6[1522];
@(posedge clk);
#1;data_in = testData6[1523];
@(posedge clk);
#1;data_in = testData6[1524];
@(posedge clk);
#1;data_in = testData6[1525];
@(posedge clk);
#1;data_in = testData6[1526];
@(posedge clk);
#1;data_in = testData6[1527];
@(posedge clk);
#1;data_in = testData6[1528];
@(posedge clk);
#1;data_in = testData6[1529];
@(posedge clk);
#1;data_in = testData6[1530];
@(posedge clk);
#1;data_in = testData6[1531];
@(posedge clk);
#1;data_in = testData6[1532];
@(posedge clk);
#1;data_in = testData6[1533];
@(posedge clk);
#1;data_in = testData6[1534];
@(posedge clk);
#1;data_in = testData6[1535];
@(posedge clk);
#1;data_in = testData6[1536];
@(posedge clk);
#1;data_in = testData6[1537];
@(posedge clk);
#1;data_in = testData6[1538];
@(posedge clk);
#1;data_in = testData6[1539];
@(posedge clk);
#1;data_in = testData6[1540];
@(posedge clk);
#1;data_in = testData6[1541];
@(posedge clk);
#1;data_in = testData6[1542];
@(posedge clk);
#1;data_in = testData6[1543];
@(posedge clk);
#1;data_in = testData6[1544];
@(posedge clk);
#1;data_in = testData6[1545];
@(posedge clk);
#1;data_in = testData6[1546];
@(posedge clk);
#1;data_in = testData6[1547];
@(posedge clk);
#1;data_in = testData6[1548];
@(posedge clk);
#1;data_in = testData6[1549];
@(posedge clk);
#1;data_in = testData6[1550];
@(posedge clk);
#1;data_in = testData6[1551];
@(posedge clk);
#1;data_in = testData6[1552];
@(posedge clk);
#1;data_in = testData6[1553];
@(posedge clk);
#1;data_in = testData6[1554];
@(posedge clk);
#1;data_in = testData6[1555];
@(posedge clk);
#1;data_in = testData6[1556];
@(posedge clk);
#1;data_in = testData6[1557];
@(posedge clk);
#1;data_in = testData6[1558];
@(posedge clk);
#1;data_in = testData6[1559];
@(posedge clk);
#1;data_in = testData6[1560];
@(posedge clk);
#1;data_in = testData6[1561];
@(posedge clk);
#1;data_in = testData6[1562];
@(posedge clk);
#1;data_in = testData6[1563];
@(posedge clk);
#1;data_in = testData6[1564];
@(posedge clk);
#1;data_in = testData6[1565];
@(posedge clk);
#1;data_in = testData6[1566];
@(posedge clk);
#1;data_in = testData6[1567];
@(posedge clk);
#1;data_in = testData6[1568];
@(posedge clk);
#1;data_in = testData6[1569];
@(posedge clk);
#1;data_in = testData6[1570];
@(posedge clk);
#1;data_in = testData6[1571];
@(posedge clk);
#1;data_in = testData6[1572];
@(posedge clk);
#1;data_in = testData6[1573];
@(posedge clk);
#1;data_in = testData6[1574];
@(posedge clk);
#1;data_in = testData6[1575];
@(posedge clk);
#1;data_in = testData6[1576];
@(posedge clk);
#1;data_in = testData6[1577];
@(posedge clk);
#1;data_in = testData6[1578];
@(posedge clk);
#1;data_in = testData6[1579];
@(posedge clk);
#1;data_in = testData6[1580];
@(posedge clk);
#1;data_in = testData6[1581];
@(posedge clk);
#1;data_in = testData6[1582];
@(posedge clk);
#1;data_in = testData6[1583];
@(posedge clk);
#1;data_in = testData6[1584];
@(posedge clk);
#1;data_in = testData6[1585];
@(posedge clk);
#1;data_in = testData6[1586];
@(posedge clk);
#1;data_in = testData6[1587];
@(posedge clk);
#1;data_in = testData6[1588];
@(posedge clk);
#1;data_in = testData6[1589];
@(posedge clk);
#1;data_in = testData6[1590];
@(posedge clk);
#1;data_in = testData6[1591];
@(posedge clk);
#1;data_in = testData6[1592];
@(posedge clk);
#1;data_in = testData6[1593];
@(posedge clk);
#1;data_in = testData6[1594];
@(posedge clk);
#1;data_in = testData6[1595];
@(posedge clk);
#1;data_in = testData6[1596];
@(posedge clk);
#1;data_in = testData6[1597];
@(posedge clk);
#1;data_in = testData6[1598];
@(posedge clk);
#1;data_in = testData6[1599];
@(posedge clk);
#1;data_in = testData6[1600];
@(posedge clk);
#1;data_in = testData6[1601];
@(posedge clk);
#1;data_in = testData6[1602];
@(posedge clk);
#1;data_in = testData6[1603];
@(posedge clk);
#1;data_in = testData6[1604];
@(posedge clk);
#1;data_in = testData6[1605];
@(posedge clk);
#1;data_in = testData6[1606];
@(posedge clk);
#1;data_in = testData6[1607];
@(posedge clk);
#1;data_in = testData6[1608];
@(posedge clk);
#1;data_in = testData6[1609];
@(posedge clk);
#1;data_in = testData6[1610];
@(posedge clk);
#1;data_in = testData6[1611];
@(posedge clk);
#1;data_in = testData6[1612];
@(posedge clk);
#1;data_in = testData6[1613];
@(posedge clk);
#1;data_in = testData6[1614];
@(posedge clk);
#1;data_in = testData6[1615];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1616]; 
@(posedge clk);
#1;data_in = testData6[1617];
@(posedge clk);
#1;data_in = testData6[1618];
@(posedge clk);
#1;data_in = testData6[1619];
@(posedge clk);
#1;data_in = testData6[1620];
@(posedge clk);
#1;data_in = testData6[1621];
@(posedge clk);
#1;data_in = testData6[1622];
@(posedge clk);
#1;data_in = testData6[1623];
@(posedge clk);
#1;data_in = testData6[1624];
@(posedge clk);
#1;data_in = testData6[1625];
@(posedge clk);
#1;data_in = testData6[1626];
@(posedge clk);
#1;data_in = testData6[1627];
@(posedge clk);
#1;data_in = testData6[1628];
@(posedge clk);
#1;data_in = testData6[1629];
@(posedge clk);
#1;data_in = testData6[1630];
@(posedge clk);
#1;data_in = testData6[1631];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1632];
@(posedge clk);
#1;data_in = testData6[1633];
@(posedge clk);
#1;data_in = testData6[1634];
@(posedge clk);
#1;data_in = testData6[1635];
@(posedge clk);
#1;data_in = testData6[1636];
@(posedge clk);
#1;data_in = testData6[1637];
@(posedge clk);
#1;data_in = testData6[1638];
@(posedge clk);
#1;data_in = testData6[1639];
@(posedge clk);
#1;data_in = testData6[1640];
@(posedge clk);
#1;data_in = testData6[1641];
@(posedge clk);
#1;data_in = testData6[1642];
@(posedge clk);
#1;data_in = testData6[1643];
@(posedge clk);
#1;data_in = testData6[1644];
@(posedge clk);
#1;data_in = testData6[1645];
@(posedge clk);
#1;data_in = testData6[1646];
@(posedge clk);
#1;data_in = testData6[1647];
@(posedge clk);
#1;data_in = testData6[1648];
@(posedge clk);
#1;data_in = testData6[1649];
@(posedge clk);
#1;data_in = testData6[1650];
@(posedge clk);
#1;data_in = testData6[1651];
@(posedge clk);
#1;data_in = testData6[1652];
@(posedge clk);
#1;data_in = testData6[1653];
@(posedge clk);
#1;data_in = testData6[1654];
@(posedge clk);
#1;data_in = testData6[1655];
@(posedge clk);
#1;data_in = testData6[1656];
@(posedge clk);
#1;data_in = testData6[1657];
@(posedge clk);
#1;data_in = testData6[1658];
@(posedge clk);
#1;data_in = testData6[1659];
@(posedge clk);
#1;data_in = testData6[1660];
@(posedge clk);
#1;data_in = testData6[1661];
@(posedge clk);
#1;data_in = testData6[1662];
@(posedge clk);
#1;data_in = testData6[1663];
@(posedge clk);
#1;data_in = testData6[1664];
@(posedge clk);
#1;data_in = testData6[1665];
@(posedge clk);
#1;data_in = testData6[1666];
@(posedge clk);
#1;data_in = testData6[1667];
@(posedge clk);
#1;data_in = testData6[1668];
@(posedge clk);
#1;data_in = testData6[1669];
@(posedge clk);
#1;data_in = testData6[1670];
@(posedge clk);
#1;data_in = testData6[1671];
@(posedge clk);
#1;data_in = testData6[1672];
@(posedge clk);
#1;data_in = testData6[1673];
@(posedge clk);
#1;data_in = testData6[1674];
@(posedge clk);
#1;data_in = testData6[1675];
@(posedge clk);
#1;data_in = testData6[1676];
@(posedge clk);
#1;data_in = testData6[1677];
@(posedge clk);
#1;data_in = testData6[1678];
@(posedge clk);
#1;data_in = testData6[1679];
@(posedge clk);
#1;data_in = testData6[1680];
@(posedge clk);
#1;data_in = testData6[1681];
@(posedge clk);
#1;data_in = testData6[1682];
@(posedge clk);
#1;data_in = testData6[1683];
@(posedge clk);
#1;data_in = testData6[1684];
@(posedge clk);
#1;data_in = testData6[1685];
@(posedge clk);
#1;data_in = testData6[1686];
@(posedge clk);
#1;data_in = testData6[1687];
@(posedge clk);
#1;data_in = testData6[1688];
@(posedge clk);
#1;data_in = testData6[1689];
@(posedge clk);
#1;data_in = testData6[1690];
@(posedge clk);
#1;data_in = testData6[1691];
@(posedge clk);
#1;data_in = testData6[1692];
@(posedge clk);
#1;data_in = testData6[1693];
@(posedge clk);
#1;data_in = testData6[1694];
@(posedge clk);
#1;data_in = testData6[1695];
@(posedge clk);
#1;data_in = testData6[1696];
@(posedge clk);
#1;data_in = testData6[1697];
@(posedge clk);
#1;data_in = testData6[1698];
@(posedge clk);
#1;data_in = testData6[1699];
@(posedge clk);
#1;data_in = testData6[1700];
@(posedge clk);
#1;data_in = testData6[1701];
@(posedge clk);
#1;data_in = testData6[1702];
@(posedge clk);
#1;data_in = testData6[1703];
@(posedge clk);
#1;data_in = testData6[1704];
@(posedge clk);
#1;data_in = testData6[1705];
@(posedge clk);
#1;data_in = testData6[1706];
@(posedge clk);
#1;data_in = testData6[1707];
@(posedge clk);
#1;data_in = testData6[1708];
@(posedge clk);
#1;data_in = testData6[1709];
@(posedge clk);
#1;data_in = testData6[1710];
@(posedge clk);
#1;data_in = testData6[1711];
@(posedge clk);
#1;data_in = testData6[1712];
@(posedge clk);
#1;data_in = testData6[1713];
@(posedge clk);
#1;data_in = testData6[1714];
@(posedge clk);
#1;data_in = testData6[1715];
@(posedge clk);
#1;data_in = testData6[1716];
@(posedge clk);
#1;data_in = testData6[1717];
@(posedge clk);
#1;data_in = testData6[1718];
@(posedge clk);
#1;data_in = testData6[1719];
@(posedge clk);
#1;data_in = testData6[1720];
@(posedge clk);
#1;data_in = testData6[1721];
@(posedge clk);
#1;data_in = testData6[1722];
@(posedge clk);
#1;data_in = testData6[1723];
@(posedge clk);
#1;data_in = testData6[1724];
@(posedge clk);
#1;data_in = testData6[1725];
@(posedge clk);
#1;data_in = testData6[1726];
@(posedge clk);
#1;data_in = testData6[1727];
@(posedge clk);
#1;data_in = testData6[1728];
@(posedge clk);
#1;data_in = testData6[1729];
@(posedge clk);
#1;data_in = testData6[1730];
@(posedge clk);
#1;data_in = testData6[1731];
@(posedge clk);
#1;data_in = testData6[1732];
@(posedge clk);
#1;data_in = testData6[1733];
@(posedge clk);
#1;data_in = testData6[1734];
@(posedge clk);
#1;data_in = testData6[1735];
@(posedge clk);
#1;data_in = testData6[1736];
@(posedge clk);
#1;data_in = testData6[1737];
@(posedge clk);
#1;data_in = testData6[1738];
@(posedge clk);
#1;data_in = testData6[1739];
@(posedge clk);
#1;data_in = testData6[1740];
@(posedge clk);
#1;data_in = testData6[1741];
@(posedge clk);
#1;data_in = testData6[1742];
@(posedge clk);
#1;data_in = testData6[1743];
@(posedge clk);
#1;data_in = testData6[1744];
@(posedge clk);
#1;data_in = testData6[1745];
@(posedge clk);
#1;data_in = testData6[1746];
@(posedge clk);
#1;data_in = testData6[1747];
@(posedge clk);
#1;data_in = testData6[1748];
@(posedge clk);
#1;data_in = testData6[1749];
@(posedge clk);
#1;data_in = testData6[1750];
@(posedge clk);
#1;data_in = testData6[1751];
@(posedge clk);
#1;data_in = testData6[1752];
@(posedge clk);
#1;data_in = testData6[1753];
@(posedge clk);
#1;data_in = testData6[1754];
@(posedge clk);
#1;data_in = testData6[1755];
@(posedge clk);
#1;data_in = testData6[1756];
@(posedge clk);
#1;data_in = testData6[1757];
@(posedge clk);
#1;data_in = testData6[1758];
@(posedge clk);
#1;data_in = testData6[1759];
@(posedge clk);
#1;data_in = testData6[1760];
@(posedge clk);
#1;data_in = testData6[1761];
@(posedge clk);
#1;data_in = testData6[1762];
@(posedge clk);
#1;data_in = testData6[1763];
@(posedge clk);
#1;data_in = testData6[1764];
@(posedge clk);
#1;data_in = testData6[1765];
@(posedge clk);
#1;data_in = testData6[1766];
@(posedge clk);
#1;data_in = testData6[1767];
@(posedge clk);
#1;data_in = testData6[1768];
@(posedge clk);
#1;data_in = testData6[1769];
@(posedge clk);
#1;data_in = testData6[1770];
@(posedge clk);
#1;data_in = testData6[1771];
@(posedge clk);
#1;data_in = testData6[1772];
@(posedge clk);
#1;data_in = testData6[1773];
@(posedge clk);
#1;data_in = testData6[1774];
@(posedge clk);
#1;data_in = testData6[1775];
@(posedge clk);
#1;data_in = testData6[1776];
@(posedge clk);
#1;data_in = testData6[1777];
@(posedge clk);
#1;data_in = testData6[1778];
@(posedge clk);
#1;data_in = testData6[1779];
@(posedge clk);
#1;data_in = testData6[1780];
@(posedge clk);
#1;data_in = testData6[1781];
@(posedge clk);
#1;data_in = testData6[1782];
@(posedge clk);
#1;data_in = testData6[1783];
@(posedge clk);
#1;data_in = testData6[1784];
@(posedge clk);
#1;data_in = testData6[1785];
@(posedge clk);
#1;data_in = testData6[1786];
@(posedge clk);
#1;data_in = testData6[1787];
@(posedge clk);
#1;data_in = testData6[1788];
@(posedge clk);
#1;data_in = testData6[1789];
@(posedge clk);
#1;data_in = testData6[1790];
@(posedge clk);
#1;data_in = testData6[1791];
@(posedge clk);
#1;data_in = testData6[1792];
@(posedge clk);
#1;data_in = testData6[1793];
@(posedge clk);
#1;data_in = testData6[1794];
@(posedge clk);
#1;data_in = testData6[1795];
@(posedge clk);
#1;data_in = testData6[1796];
@(posedge clk);
#1;data_in = testData6[1797];
@(posedge clk);
#1;data_in = testData6[1798];
@(posedge clk);
#1;data_in = testData6[1799];
@(posedge clk);
#1;data_in = testData6[1800];
@(posedge clk);
#1;data_in = testData6[1801];
@(posedge clk);
#1;data_in = testData6[1802];
@(posedge clk);
#1;data_in = testData6[1803];
@(posedge clk);
#1;data_in = testData6[1804];
@(posedge clk);
#1;data_in = testData6[1805];
@(posedge clk);
#1;data_in = testData6[1806];
@(posedge clk);
#1;data_in = testData6[1807];
@(posedge clk);
#1;data_in = testData6[1808];
@(posedge clk);
#1;data_in = testData6[1809];
@(posedge clk);
#1;data_in = testData6[1810];
@(posedge clk);
#1;data_in = testData6[1811];
@(posedge clk);
#1;data_in = testData6[1812];
@(posedge clk);
#1;data_in = testData6[1813];
@(posedge clk);
#1;data_in = testData6[1814];
@(posedge clk);
#1;data_in = testData6[1815];
@(posedge clk);
#1;data_in = testData6[1816];
@(posedge clk);
#1;data_in = testData6[1817];
@(posedge clk);
#1;data_in = testData6[1818];
@(posedge clk);
#1;data_in = testData6[1819];
@(posedge clk);
#1;data_in = testData6[1820];
@(posedge clk);
#1;data_in = testData6[1821];
@(posedge clk);
#1;data_in = testData6[1822];
@(posedge clk);
#1;data_in = testData6[1823];
@(posedge clk);
#1;data_in = testData6[1824];
@(posedge clk);
#1;data_in = testData6[1825];
@(posedge clk);
#1;data_in = testData6[1826];
@(posedge clk);
#1;data_in = testData6[1827];
@(posedge clk);
#1;data_in = testData6[1828];
@(posedge clk);
#1;data_in = testData6[1829];
@(posedge clk);
#1;data_in = testData6[1830];
@(posedge clk);
#1;data_in = testData6[1831];
@(posedge clk);
#1;data_in = testData6[1832];
@(posedge clk);
#1;data_in = testData6[1833];
@(posedge clk);
#1;data_in = testData6[1834];
@(posedge clk);
#1;data_in = testData6[1835];
@(posedge clk);
#1;data_in = testData6[1836];
@(posedge clk);
#1;data_in = testData6[1837];
@(posedge clk);
#1;data_in = testData6[1838];
@(posedge clk);
#1;data_in = testData6[1839];
@(posedge clk);
#1;data_in = testData6[1840];
@(posedge clk);
#1;data_in = testData6[1841];
@(posedge clk);
#1;data_in = testData6[1842];
@(posedge clk);
#1;data_in = testData6[1843];
@(posedge clk);
#1;data_in = testData6[1844];
@(posedge clk);
#1;data_in = testData6[1845];
@(posedge clk);
#1;data_in = testData6[1846];
@(posedge clk);
#1;data_in = testData6[1847];
@(posedge clk);
#1;data_in = testData6[1848];
@(posedge clk);
#1;data_in = testData6[1849];
@(posedge clk);
#1;data_in = testData6[1850];
@(posedge clk);
#1;data_in = testData6[1851];
@(posedge clk);
#1;data_in = testData6[1852];
@(posedge clk);
#1;data_in = testData6[1853];
@(posedge clk);
#1;data_in = testData6[1854];
@(posedge clk);
#1;data_in = testData6[1855];
@(posedge clk);
#1;data_in = testData6[1856];
@(posedge clk);
#1;data_in = testData6[1857];
@(posedge clk);
#1;data_in = testData6[1858];
@(posedge clk);
#1;data_in = testData6[1859];
@(posedge clk);
#1;data_in = testData6[1860];
@(posedge clk);
#1;data_in = testData6[1861];
@(posedge clk);
#1;data_in = testData6[1862];
@(posedge clk);
#1;data_in = testData6[1863];
@(posedge clk);
#1;data_in = testData6[1864];
@(posedge clk);
#1;data_in = testData6[1865];
@(posedge clk);
#1;data_in = testData6[1866];
@(posedge clk);
#1;data_in = testData6[1867];
@(posedge clk);
#1;data_in = testData6[1868];
@(posedge clk);
#1;data_in = testData6[1869];
@(posedge clk);
#1;data_in = testData6[1870];
@(posedge clk);
#1;data_in = testData6[1871];
@(posedge clk);
#1;data_in = testData6[1872];
@(posedge clk);
#1;data_in = testData6[1873];
@(posedge clk);
#1;data_in = testData6[1874];
@(posedge clk);
#1;data_in = testData6[1875];
@(posedge clk);
#1;data_in = testData6[1876];
@(posedge clk);
#1;data_in = testData6[1877];
@(posedge clk);
#1;data_in = testData6[1878];
@(posedge clk);
#1;data_in = testData6[1879];
@(posedge clk);
#1;data_in = testData6[1880];
@(posedge clk);
#1;data_in = testData6[1881];
@(posedge clk);
#1;data_in = testData6[1882];
@(posedge clk);
#1;data_in = testData6[1883];
@(posedge clk);
#1;data_in = testData6[1884];
@(posedge clk);
#1;data_in = testData6[1885];
@(posedge clk);
#1;data_in = testData6[1886];
@(posedge clk);
#1;data_in = testData6[1887];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1888]; 
@(posedge clk);
#1;data_in = testData6[1889];
@(posedge clk);
#1;data_in = testData6[1890];
@(posedge clk);
#1;data_in = testData6[1891];
@(posedge clk);
#1;data_in = testData6[1892];
@(posedge clk);
#1;data_in = testData6[1893];
@(posedge clk);
#1;data_in = testData6[1894];
@(posedge clk);
#1;data_in = testData6[1895];
@(posedge clk);
#1;data_in = testData6[1896];
@(posedge clk);
#1;data_in = testData6[1897];
@(posedge clk);
#1;data_in = testData6[1898];
@(posedge clk);
#1;data_in = testData6[1899];
@(posedge clk);
#1;data_in = testData6[1900];
@(posedge clk);
#1;data_in = testData6[1901];
@(posedge clk);
#1;data_in = testData6[1902];
@(posedge clk);
#1;data_in = testData6[1903];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1904];
@(posedge clk);
#1;data_in = testData6[1905];
@(posedge clk);
#1;data_in = testData6[1906];
@(posedge clk);
#1;data_in = testData6[1907];
@(posedge clk);
#1;data_in = testData6[1908];
@(posedge clk);
#1;data_in = testData6[1909];
@(posedge clk);
#1;data_in = testData6[1910];
@(posedge clk);
#1;data_in = testData6[1911];
@(posedge clk);
#1;data_in = testData6[1912];
@(posedge clk);
#1;data_in = testData6[1913];
@(posedge clk);
#1;data_in = testData6[1914];
@(posedge clk);
#1;data_in = testData6[1915];
@(posedge clk);
#1;data_in = testData6[1916];
@(posedge clk);
#1;data_in = testData6[1917];
@(posedge clk);
#1;data_in = testData6[1918];
@(posedge clk);
#1;data_in = testData6[1919];
@(posedge clk);
#1;data_in = testData6[1920];
@(posedge clk);
#1;data_in = testData6[1921];
@(posedge clk);
#1;data_in = testData6[1922];
@(posedge clk);
#1;data_in = testData6[1923];
@(posedge clk);
#1;data_in = testData6[1924];
@(posedge clk);
#1;data_in = testData6[1925];
@(posedge clk);
#1;data_in = testData6[1926];
@(posedge clk);
#1;data_in = testData6[1927];
@(posedge clk);
#1;data_in = testData6[1928];
@(posedge clk);
#1;data_in = testData6[1929];
@(posedge clk);
#1;data_in = testData6[1930];
@(posedge clk);
#1;data_in = testData6[1931];
@(posedge clk);
#1;data_in = testData6[1932];
@(posedge clk);
#1;data_in = testData6[1933];
@(posedge clk);
#1;data_in = testData6[1934];
@(posedge clk);
#1;data_in = testData6[1935];
@(posedge clk);
#1;data_in = testData6[1936];
@(posedge clk);
#1;data_in = testData6[1937];
@(posedge clk);
#1;data_in = testData6[1938];
@(posedge clk);
#1;data_in = testData6[1939];
@(posedge clk);
#1;data_in = testData6[1940];
@(posedge clk);
#1;data_in = testData6[1941];
@(posedge clk);
#1;data_in = testData6[1942];
@(posedge clk);
#1;data_in = testData6[1943];
@(posedge clk);
#1;data_in = testData6[1944];
@(posedge clk);
#1;data_in = testData6[1945];
@(posedge clk);
#1;data_in = testData6[1946];
@(posedge clk);
#1;data_in = testData6[1947];
@(posedge clk);
#1;data_in = testData6[1948];
@(posedge clk);
#1;data_in = testData6[1949];
@(posedge clk);
#1;data_in = testData6[1950];
@(posedge clk);
#1;data_in = testData6[1951];
@(posedge clk);
#1;data_in = testData6[1952];
@(posedge clk);
#1;data_in = testData6[1953];
@(posedge clk);
#1;data_in = testData6[1954];
@(posedge clk);
#1;data_in = testData6[1955];
@(posedge clk);
#1;data_in = testData6[1956];
@(posedge clk);
#1;data_in = testData6[1957];
@(posedge clk);
#1;data_in = testData6[1958];
@(posedge clk);
#1;data_in = testData6[1959];
@(posedge clk);
#1;data_in = testData6[1960];
@(posedge clk);
#1;data_in = testData6[1961];
@(posedge clk);
#1;data_in = testData6[1962];
@(posedge clk);
#1;data_in = testData6[1963];
@(posedge clk);
#1;data_in = testData6[1964];
@(posedge clk);
#1;data_in = testData6[1965];
@(posedge clk);
#1;data_in = testData6[1966];
@(posedge clk);
#1;data_in = testData6[1967];
@(posedge clk);
#1;data_in = testData6[1968];
@(posedge clk);
#1;data_in = testData6[1969];
@(posedge clk);
#1;data_in = testData6[1970];
@(posedge clk);
#1;data_in = testData6[1971];
@(posedge clk);
#1;data_in = testData6[1972];
@(posedge clk);
#1;data_in = testData6[1973];
@(posedge clk);
#1;data_in = testData6[1974];
@(posedge clk);
#1;data_in = testData6[1975];
@(posedge clk);
#1;data_in = testData6[1976];
@(posedge clk);
#1;data_in = testData6[1977];
@(posedge clk);
#1;data_in = testData6[1978];
@(posedge clk);
#1;data_in = testData6[1979];
@(posedge clk);
#1;data_in = testData6[1980];
@(posedge clk);
#1;data_in = testData6[1981];
@(posedge clk);
#1;data_in = testData6[1982];
@(posedge clk);
#1;data_in = testData6[1983];
@(posedge clk);
#1;data_in = testData6[1984];
@(posedge clk);
#1;data_in = testData6[1985];
@(posedge clk);
#1;data_in = testData6[1986];
@(posedge clk);
#1;data_in = testData6[1987];
@(posedge clk);
#1;data_in = testData6[1988];
@(posedge clk);
#1;data_in = testData6[1989];
@(posedge clk);
#1;data_in = testData6[1990];
@(posedge clk);
#1;data_in = testData6[1991];
@(posedge clk);
#1;data_in = testData6[1992];
@(posedge clk);
#1;data_in = testData6[1993];
@(posedge clk);
#1;data_in = testData6[1994];
@(posedge clk);
#1;data_in = testData6[1995];
@(posedge clk);
#1;data_in = testData6[1996];
@(posedge clk);
#1;data_in = testData6[1997];
@(posedge clk);
#1;data_in = testData6[1998];
@(posedge clk);
#1;data_in = testData6[1999];
@(posedge clk);
#1;data_in = testData6[2000];
@(posedge clk);
#1;data_in = testData6[2001];
@(posedge clk);
#1;data_in = testData6[2002];
@(posedge clk);
#1;data_in = testData6[2003];
@(posedge clk);
#1;data_in = testData6[2004];
@(posedge clk);
#1;data_in = testData6[2005];
@(posedge clk);
#1;data_in = testData6[2006];
@(posedge clk);
#1;data_in = testData6[2007];
@(posedge clk);
#1;data_in = testData6[2008];
@(posedge clk);
#1;data_in = testData6[2009];
@(posedge clk);
#1;data_in = testData6[2010];
@(posedge clk);
#1;data_in = testData6[2011];
@(posedge clk);
#1;data_in = testData6[2012];
@(posedge clk);
#1;data_in = testData6[2013];
@(posedge clk);
#1;data_in = testData6[2014];
@(posedge clk);
#1;data_in = testData6[2015];
@(posedge clk);
#1;data_in = testData6[2016];
@(posedge clk);
#1;data_in = testData6[2017];
@(posedge clk);
#1;data_in = testData6[2018];
@(posedge clk);
#1;data_in = testData6[2019];
@(posedge clk);
#1;data_in = testData6[2020];
@(posedge clk);
#1;data_in = testData6[2021];
@(posedge clk);
#1;data_in = testData6[2022];
@(posedge clk);
#1;data_in = testData6[2023];
@(posedge clk);
#1;data_in = testData6[2024];
@(posedge clk);
#1;data_in = testData6[2025];
@(posedge clk);
#1;data_in = testData6[2026];
@(posedge clk);
#1;data_in = testData6[2027];
@(posedge clk);
#1;data_in = testData6[2028];
@(posedge clk);
#1;data_in = testData6[2029];
@(posedge clk);
#1;data_in = testData6[2030];
@(posedge clk);
#1;data_in = testData6[2031];
@(posedge clk);
#1;data_in = testData6[2032];
@(posedge clk);
#1;data_in = testData6[2033];
@(posedge clk);
#1;data_in = testData6[2034];
@(posedge clk);
#1;data_in = testData6[2035];
@(posedge clk);
#1;data_in = testData6[2036];
@(posedge clk);
#1;data_in = testData6[2037];
@(posedge clk);
#1;data_in = testData6[2038];
@(posedge clk);
#1;data_in = testData6[2039];
@(posedge clk);
#1;data_in = testData6[2040];
@(posedge clk);
#1;data_in = testData6[2041];
@(posedge clk);
#1;data_in = testData6[2042];
@(posedge clk);
#1;data_in = testData6[2043];
@(posedge clk);
#1;data_in = testData6[2044];
@(posedge clk);
#1;data_in = testData6[2045];
@(posedge clk);
#1;data_in = testData6[2046];
@(posedge clk);
#1;data_in = testData6[2047];
@(posedge clk);
#1;data_in = testData6[2048];
@(posedge clk);
#1;data_in = testData6[2049];
@(posedge clk);
#1;data_in = testData6[2050];
@(posedge clk);
#1;data_in = testData6[2051];
@(posedge clk);
#1;data_in = testData6[2052];
@(posedge clk);
#1;data_in = testData6[2053];
@(posedge clk);
#1;data_in = testData6[2054];
@(posedge clk);
#1;data_in = testData6[2055];
@(posedge clk);
#1;data_in = testData6[2056];
@(posedge clk);
#1;data_in = testData6[2057];
@(posedge clk);
#1;data_in = testData6[2058];
@(posedge clk);
#1;data_in = testData6[2059];
@(posedge clk);
#1;data_in = testData6[2060];
@(posedge clk);
#1;data_in = testData6[2061];
@(posedge clk);
#1;data_in = testData6[2062];
@(posedge clk);
#1;data_in = testData6[2063];
@(posedge clk);
#1;data_in = testData6[2064];
@(posedge clk);
#1;data_in = testData6[2065];
@(posedge clk);
#1;data_in = testData6[2066];
@(posedge clk);
#1;data_in = testData6[2067];
@(posedge clk);
#1;data_in = testData6[2068];
@(posedge clk);
#1;data_in = testData6[2069];
@(posedge clk);
#1;data_in = testData6[2070];
@(posedge clk);
#1;data_in = testData6[2071];
@(posedge clk);
#1;data_in = testData6[2072];
@(posedge clk);
#1;data_in = testData6[2073];
@(posedge clk);
#1;data_in = testData6[2074];
@(posedge clk);
#1;data_in = testData6[2075];
@(posedge clk);
#1;data_in = testData6[2076];
@(posedge clk);
#1;data_in = testData6[2077];
@(posedge clk);
#1;data_in = testData6[2078];
@(posedge clk);
#1;data_in = testData6[2079];
@(posedge clk);
#1;data_in = testData6[2080];
@(posedge clk);
#1;data_in = testData6[2081];
@(posedge clk);
#1;data_in = testData6[2082];
@(posedge clk);
#1;data_in = testData6[2083];
@(posedge clk);
#1;data_in = testData6[2084];
@(posedge clk);
#1;data_in = testData6[2085];
@(posedge clk);
#1;data_in = testData6[2086];
@(posedge clk);
#1;data_in = testData6[2087];
@(posedge clk);
#1;data_in = testData6[2088];
@(posedge clk);
#1;data_in = testData6[2089];
@(posedge clk);
#1;data_in = testData6[2090];
@(posedge clk);
#1;data_in = testData6[2091];
@(posedge clk);
#1;data_in = testData6[2092];
@(posedge clk);
#1;data_in = testData6[2093];
@(posedge clk);
#1;data_in = testData6[2094];
@(posedge clk);
#1;data_in = testData6[2095];
@(posedge clk);
#1;data_in = testData6[2096];
@(posedge clk);
#1;data_in = testData6[2097];
@(posedge clk);
#1;data_in = testData6[2098];
@(posedge clk);
#1;data_in = testData6[2099];
@(posedge clk);
#1;data_in = testData6[2100];
@(posedge clk);
#1;data_in = testData6[2101];
@(posedge clk);
#1;data_in = testData6[2102];
@(posedge clk);
#1;data_in = testData6[2103];
@(posedge clk);
#1;data_in = testData6[2104];
@(posedge clk);
#1;data_in = testData6[2105];
@(posedge clk);
#1;data_in = testData6[2106];
@(posedge clk);
#1;data_in = testData6[2107];
@(posedge clk);
#1;data_in = testData6[2108];
@(posedge clk);
#1;data_in = testData6[2109];
@(posedge clk);
#1;data_in = testData6[2110];
@(posedge clk);
#1;data_in = testData6[2111];
@(posedge clk);
#1;data_in = testData6[2112];
@(posedge clk);
#1;data_in = testData6[2113];
@(posedge clk);
#1;data_in = testData6[2114];
@(posedge clk);
#1;data_in = testData6[2115];
@(posedge clk);
#1;data_in = testData6[2116];
@(posedge clk);
#1;data_in = testData6[2117];
@(posedge clk);
#1;data_in = testData6[2118];
@(posedge clk);
#1;data_in = testData6[2119];
@(posedge clk);
#1;data_in = testData6[2120];
@(posedge clk);
#1;data_in = testData6[2121];
@(posedge clk);
#1;data_in = testData6[2122];
@(posedge clk);
#1;data_in = testData6[2123];
@(posedge clk);
#1;data_in = testData6[2124];
@(posedge clk);
#1;data_in = testData6[2125];
@(posedge clk);
#1;data_in = testData6[2126];
@(posedge clk);
#1;data_in = testData6[2127];
@(posedge clk);
#1;data_in = testData6[2128];
@(posedge clk);
#1;data_in = testData6[2129];
@(posedge clk);
#1;data_in = testData6[2130];
@(posedge clk);
#1;data_in = testData6[2131];
@(posedge clk);
#1;data_in = testData6[2132];
@(posedge clk);
#1;data_in = testData6[2133];
@(posedge clk);
#1;data_in = testData6[2134];
@(posedge clk);
#1;data_in = testData6[2135];
@(posedge clk);
#1;data_in = testData6[2136];
@(posedge clk);
#1;data_in = testData6[2137];
@(posedge clk);
#1;data_in = testData6[2138];
@(posedge clk);
#1;data_in = testData6[2139];
@(posedge clk);
#1;data_in = testData6[2140];
@(posedge clk);
#1;data_in = testData6[2141];
@(posedge clk);
#1;data_in = testData6[2142];
@(posedge clk);
#1;data_in = testData6[2143];
@(posedge clk);
#1;data_in = testData6[2144];
@(posedge clk);
#1;data_in = testData6[2145];
@(posedge clk);
#1;data_in = testData6[2146];
@(posedge clk);
#1;data_in = testData6[2147];
@(posedge clk);
#1;data_in = testData6[2148];
@(posedge clk);
#1;data_in = testData6[2149];
@(posedge clk);
#1;data_in = testData6[2150];
@(posedge clk);
#1;data_in = testData6[2151];
@(posedge clk);
#1;data_in = testData6[2152];
@(posedge clk);
#1;data_in = testData6[2153];
@(posedge clk);
#1;data_in = testData6[2154];
@(posedge clk);
#1;data_in = testData6[2155];
@(posedge clk);
#1;data_in = testData6[2156];
@(posedge clk);
#1;data_in = testData6[2157];
@(posedge clk);
#1;data_in = testData6[2158];
@(posedge clk);
#1;data_in = testData6[2159];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2160]; 
@(posedge clk);
#1;data_in = testData6[2161];
@(posedge clk);
#1;data_in = testData6[2162];
@(posedge clk);
#1;data_in = testData6[2163];
@(posedge clk);
#1;data_in = testData6[2164];
@(posedge clk);
#1;data_in = testData6[2165];
@(posedge clk);
#1;data_in = testData6[2166];
@(posedge clk);
#1;data_in = testData6[2167];
@(posedge clk);
#1;data_in = testData6[2168];
@(posedge clk);
#1;data_in = testData6[2169];
@(posedge clk);
#1;data_in = testData6[2170];
@(posedge clk);
#1;data_in = testData6[2171];
@(posedge clk);
#1;data_in = testData6[2172];
@(posedge clk);
#1;data_in = testData6[2173];
@(posedge clk);
#1;data_in = testData6[2174];
@(posedge clk);
#1;data_in = testData6[2175];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2176];
@(posedge clk);
#1;data_in = testData6[2177];
@(posedge clk);
#1;data_in = testData6[2178];
@(posedge clk);
#1;data_in = testData6[2179];
@(posedge clk);
#1;data_in = testData6[2180];
@(posedge clk);
#1;data_in = testData6[2181];
@(posedge clk);
#1;data_in = testData6[2182];
@(posedge clk);
#1;data_in = testData6[2183];
@(posedge clk);
#1;data_in = testData6[2184];
@(posedge clk);
#1;data_in = testData6[2185];
@(posedge clk);
#1;data_in = testData6[2186];
@(posedge clk);
#1;data_in = testData6[2187];
@(posedge clk);
#1;data_in = testData6[2188];
@(posedge clk);
#1;data_in = testData6[2189];
@(posedge clk);
#1;data_in = testData6[2190];
@(posedge clk);
#1;data_in = testData6[2191];
@(posedge clk);
#1;data_in = testData6[2192];
@(posedge clk);
#1;data_in = testData6[2193];
@(posedge clk);
#1;data_in = testData6[2194];
@(posedge clk);
#1;data_in = testData6[2195];
@(posedge clk);
#1;data_in = testData6[2196];
@(posedge clk);
#1;data_in = testData6[2197];
@(posedge clk);
#1;data_in = testData6[2198];
@(posedge clk);
#1;data_in = testData6[2199];
@(posedge clk);
#1;data_in = testData6[2200];
@(posedge clk);
#1;data_in = testData6[2201];
@(posedge clk);
#1;data_in = testData6[2202];
@(posedge clk);
#1;data_in = testData6[2203];
@(posedge clk);
#1;data_in = testData6[2204];
@(posedge clk);
#1;data_in = testData6[2205];
@(posedge clk);
#1;data_in = testData6[2206];
@(posedge clk);
#1;data_in = testData6[2207];
@(posedge clk);
#1;data_in = testData6[2208];
@(posedge clk);
#1;data_in = testData6[2209];
@(posedge clk);
#1;data_in = testData6[2210];
@(posedge clk);
#1;data_in = testData6[2211];
@(posedge clk);
#1;data_in = testData6[2212];
@(posedge clk);
#1;data_in = testData6[2213];
@(posedge clk);
#1;data_in = testData6[2214];
@(posedge clk);
#1;data_in = testData6[2215];
@(posedge clk);
#1;data_in = testData6[2216];
@(posedge clk);
#1;data_in = testData6[2217];
@(posedge clk);
#1;data_in = testData6[2218];
@(posedge clk);
#1;data_in = testData6[2219];
@(posedge clk);
#1;data_in = testData6[2220];
@(posedge clk);
#1;data_in = testData6[2221];
@(posedge clk);
#1;data_in = testData6[2222];
@(posedge clk);
#1;data_in = testData6[2223];
@(posedge clk);
#1;data_in = testData6[2224];
@(posedge clk);
#1;data_in = testData6[2225];
@(posedge clk);
#1;data_in = testData6[2226];
@(posedge clk);
#1;data_in = testData6[2227];
@(posedge clk);
#1;data_in = testData6[2228];
@(posedge clk);
#1;data_in = testData6[2229];
@(posedge clk);
#1;data_in = testData6[2230];
@(posedge clk);
#1;data_in = testData6[2231];
@(posedge clk);
#1;data_in = testData6[2232];
@(posedge clk);
#1;data_in = testData6[2233];
@(posedge clk);
#1;data_in = testData6[2234];
@(posedge clk);
#1;data_in = testData6[2235];
@(posedge clk);
#1;data_in = testData6[2236];
@(posedge clk);
#1;data_in = testData6[2237];
@(posedge clk);
#1;data_in = testData6[2238];
@(posedge clk);
#1;data_in = testData6[2239];
@(posedge clk);
#1;data_in = testData6[2240];
@(posedge clk);
#1;data_in = testData6[2241];
@(posedge clk);
#1;data_in = testData6[2242];
@(posedge clk);
#1;data_in = testData6[2243];
@(posedge clk);
#1;data_in = testData6[2244];
@(posedge clk);
#1;data_in = testData6[2245];
@(posedge clk);
#1;data_in = testData6[2246];
@(posedge clk);
#1;data_in = testData6[2247];
@(posedge clk);
#1;data_in = testData6[2248];
@(posedge clk);
#1;data_in = testData6[2249];
@(posedge clk);
#1;data_in = testData6[2250];
@(posedge clk);
#1;data_in = testData6[2251];
@(posedge clk);
#1;data_in = testData6[2252];
@(posedge clk);
#1;data_in = testData6[2253];
@(posedge clk);
#1;data_in = testData6[2254];
@(posedge clk);
#1;data_in = testData6[2255];
@(posedge clk);
#1;data_in = testData6[2256];
@(posedge clk);
#1;data_in = testData6[2257];
@(posedge clk);
#1;data_in = testData6[2258];
@(posedge clk);
#1;data_in = testData6[2259];
@(posedge clk);
#1;data_in = testData6[2260];
@(posedge clk);
#1;data_in = testData6[2261];
@(posedge clk);
#1;data_in = testData6[2262];
@(posedge clk);
#1;data_in = testData6[2263];
@(posedge clk);
#1;data_in = testData6[2264];
@(posedge clk);
#1;data_in = testData6[2265];
@(posedge clk);
#1;data_in = testData6[2266];
@(posedge clk);
#1;data_in = testData6[2267];
@(posedge clk);
#1;data_in = testData6[2268];
@(posedge clk);
#1;data_in = testData6[2269];
@(posedge clk);
#1;data_in = testData6[2270];
@(posedge clk);
#1;data_in = testData6[2271];
@(posedge clk);
#1;data_in = testData6[2272];
@(posedge clk);
#1;data_in = testData6[2273];
@(posedge clk);
#1;data_in = testData6[2274];
@(posedge clk);
#1;data_in = testData6[2275];
@(posedge clk);
#1;data_in = testData6[2276];
@(posedge clk);
#1;data_in = testData6[2277];
@(posedge clk);
#1;data_in = testData6[2278];
@(posedge clk);
#1;data_in = testData6[2279];
@(posedge clk);
#1;data_in = testData6[2280];
@(posedge clk);
#1;data_in = testData6[2281];
@(posedge clk);
#1;data_in = testData6[2282];
@(posedge clk);
#1;data_in = testData6[2283];
@(posedge clk);
#1;data_in = testData6[2284];
@(posedge clk);
#1;data_in = testData6[2285];
@(posedge clk);
#1;data_in = testData6[2286];
@(posedge clk);
#1;data_in = testData6[2287];
@(posedge clk);
#1;data_in = testData6[2288];
@(posedge clk);
#1;data_in = testData6[2289];
@(posedge clk);
#1;data_in = testData6[2290];
@(posedge clk);
#1;data_in = testData6[2291];
@(posedge clk);
#1;data_in = testData6[2292];
@(posedge clk);
#1;data_in = testData6[2293];
@(posedge clk);
#1;data_in = testData6[2294];
@(posedge clk);
#1;data_in = testData6[2295];
@(posedge clk);
#1;data_in = testData6[2296];
@(posedge clk);
#1;data_in = testData6[2297];
@(posedge clk);
#1;data_in = testData6[2298];
@(posedge clk);
#1;data_in = testData6[2299];
@(posedge clk);
#1;data_in = testData6[2300];
@(posedge clk);
#1;data_in = testData6[2301];
@(posedge clk);
#1;data_in = testData6[2302];
@(posedge clk);
#1;data_in = testData6[2303];
@(posedge clk);
#1;data_in = testData6[2304];
@(posedge clk);
#1;data_in = testData6[2305];
@(posedge clk);
#1;data_in = testData6[2306];
@(posedge clk);
#1;data_in = testData6[2307];
@(posedge clk);
#1;data_in = testData6[2308];
@(posedge clk);
#1;data_in = testData6[2309];
@(posedge clk);
#1;data_in = testData6[2310];
@(posedge clk);
#1;data_in = testData6[2311];
@(posedge clk);
#1;data_in = testData6[2312];
@(posedge clk);
#1;data_in = testData6[2313];
@(posedge clk);
#1;data_in = testData6[2314];
@(posedge clk);
#1;data_in = testData6[2315];
@(posedge clk);
#1;data_in = testData6[2316];
@(posedge clk);
#1;data_in = testData6[2317];
@(posedge clk);
#1;data_in = testData6[2318];
@(posedge clk);
#1;data_in = testData6[2319];
@(posedge clk);
#1;data_in = testData6[2320];
@(posedge clk);
#1;data_in = testData6[2321];
@(posedge clk);
#1;data_in = testData6[2322];
@(posedge clk);
#1;data_in = testData6[2323];
@(posedge clk);
#1;data_in = testData6[2324];
@(posedge clk);
#1;data_in = testData6[2325];
@(posedge clk);
#1;data_in = testData6[2326];
@(posedge clk);
#1;data_in = testData6[2327];
@(posedge clk);
#1;data_in = testData6[2328];
@(posedge clk);
#1;data_in = testData6[2329];
@(posedge clk);
#1;data_in = testData6[2330];
@(posedge clk);
#1;data_in = testData6[2331];
@(posedge clk);
#1;data_in = testData6[2332];
@(posedge clk);
#1;data_in = testData6[2333];
@(posedge clk);
#1;data_in = testData6[2334];
@(posedge clk);
#1;data_in = testData6[2335];
@(posedge clk);
#1;data_in = testData6[2336];
@(posedge clk);
#1;data_in = testData6[2337];
@(posedge clk);
#1;data_in = testData6[2338];
@(posedge clk);
#1;data_in = testData6[2339];
@(posedge clk);
#1;data_in = testData6[2340];
@(posedge clk);
#1;data_in = testData6[2341];
@(posedge clk);
#1;data_in = testData6[2342];
@(posedge clk);
#1;data_in = testData6[2343];
@(posedge clk);
#1;data_in = testData6[2344];
@(posedge clk);
#1;data_in = testData6[2345];
@(posedge clk);
#1;data_in = testData6[2346];
@(posedge clk);
#1;data_in = testData6[2347];
@(posedge clk);
#1;data_in = testData6[2348];
@(posedge clk);
#1;data_in = testData6[2349];
@(posedge clk);
#1;data_in = testData6[2350];
@(posedge clk);
#1;data_in = testData6[2351];
@(posedge clk);
#1;data_in = testData6[2352];
@(posedge clk);
#1;data_in = testData6[2353];
@(posedge clk);
#1;data_in = testData6[2354];
@(posedge clk);
#1;data_in = testData6[2355];
@(posedge clk);
#1;data_in = testData6[2356];
@(posedge clk);
#1;data_in = testData6[2357];
@(posedge clk);
#1;data_in = testData6[2358];
@(posedge clk);
#1;data_in = testData6[2359];
@(posedge clk);
#1;data_in = testData6[2360];
@(posedge clk);
#1;data_in = testData6[2361];
@(posedge clk);
#1;data_in = testData6[2362];
@(posedge clk);
#1;data_in = testData6[2363];
@(posedge clk);
#1;data_in = testData6[2364];
@(posedge clk);
#1;data_in = testData6[2365];
@(posedge clk);
#1;data_in = testData6[2366];
@(posedge clk);
#1;data_in = testData6[2367];
@(posedge clk);
#1;data_in = testData6[2368];
@(posedge clk);
#1;data_in = testData6[2369];
@(posedge clk);
#1;data_in = testData6[2370];
@(posedge clk);
#1;data_in = testData6[2371];
@(posedge clk);
#1;data_in = testData6[2372];
@(posedge clk);
#1;data_in = testData6[2373];
@(posedge clk);
#1;data_in = testData6[2374];
@(posedge clk);
#1;data_in = testData6[2375];
@(posedge clk);
#1;data_in = testData6[2376];
@(posedge clk);
#1;data_in = testData6[2377];
@(posedge clk);
#1;data_in = testData6[2378];
@(posedge clk);
#1;data_in = testData6[2379];
@(posedge clk);
#1;data_in = testData6[2380];
@(posedge clk);
#1;data_in = testData6[2381];
@(posedge clk);
#1;data_in = testData6[2382];
@(posedge clk);
#1;data_in = testData6[2383];
@(posedge clk);
#1;data_in = testData6[2384];
@(posedge clk);
#1;data_in = testData6[2385];
@(posedge clk);
#1;data_in = testData6[2386];
@(posedge clk);
#1;data_in = testData6[2387];
@(posedge clk);
#1;data_in = testData6[2388];
@(posedge clk);
#1;data_in = testData6[2389];
@(posedge clk);
#1;data_in = testData6[2390];
@(posedge clk);
#1;data_in = testData6[2391];
@(posedge clk);
#1;data_in = testData6[2392];
@(posedge clk);
#1;data_in = testData6[2393];
@(posedge clk);
#1;data_in = testData6[2394];
@(posedge clk);
#1;data_in = testData6[2395];
@(posedge clk);
#1;data_in = testData6[2396];
@(posedge clk);
#1;data_in = testData6[2397];
@(posedge clk);
#1;data_in = testData6[2398];
@(posedge clk);
#1;data_in = testData6[2399];
@(posedge clk);
#1;data_in = testData6[2400];
@(posedge clk);
#1;data_in = testData6[2401];
@(posedge clk);
#1;data_in = testData6[2402];
@(posedge clk);
#1;data_in = testData6[2403];
@(posedge clk);
#1;data_in = testData6[2404];
@(posedge clk);
#1;data_in = testData6[2405];
@(posedge clk);
#1;data_in = testData6[2406];
@(posedge clk);
#1;data_in = testData6[2407];
@(posedge clk);
#1;data_in = testData6[2408];
@(posedge clk);
#1;data_in = testData6[2409];
@(posedge clk);
#1;data_in = testData6[2410];
@(posedge clk);
#1;data_in = testData6[2411];
@(posedge clk);
#1;data_in = testData6[2412];
@(posedge clk);
#1;data_in = testData6[2413];
@(posedge clk);
#1;data_in = testData6[2414];
@(posedge clk);
#1;data_in = testData6[2415];
@(posedge clk);
#1;data_in = testData6[2416];
@(posedge clk);
#1;data_in = testData6[2417];
@(posedge clk);
#1;data_in = testData6[2418];
@(posedge clk);
#1;data_in = testData6[2419];
@(posedge clk);
#1;data_in = testData6[2420];
@(posedge clk);
#1;data_in = testData6[2421];
@(posedge clk);
#1;data_in = testData6[2422];
@(posedge clk);
#1;data_in = testData6[2423];
@(posedge clk);
#1;data_in = testData6[2424];
@(posedge clk);
#1;data_in = testData6[2425];
@(posedge clk);
#1;data_in = testData6[2426];
@(posedge clk);
#1;data_in = testData6[2427];
@(posedge clk);
#1;data_in = testData6[2428];
@(posedge clk);
#1;data_in = testData6[2429];
@(posedge clk);
#1;data_in = testData6[2430];
@(posedge clk);
#1;data_in = testData6[2431];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2432]; 
@(posedge clk);
#1;data_in = testData6[2433];
@(posedge clk);
#1;data_in = testData6[2434];
@(posedge clk);
#1;data_in = testData6[2435];
@(posedge clk);
#1;data_in = testData6[2436];
@(posedge clk);
#1;data_in = testData6[2437];
@(posedge clk);
#1;data_in = testData6[2438];
@(posedge clk);
#1;data_in = testData6[2439];
@(posedge clk);
#1;data_in = testData6[2440];
@(posedge clk);
#1;data_in = testData6[2441];
@(posedge clk);
#1;data_in = testData6[2442];
@(posedge clk);
#1;data_in = testData6[2443];
@(posedge clk);
#1;data_in = testData6[2444];
@(posedge clk);
#1;data_in = testData6[2445];
@(posedge clk);
#1;data_in = testData6[2446];
@(posedge clk);
#1;data_in = testData6[2447];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2448];
@(posedge clk);
#1;data_in = testData6[2449];
@(posedge clk);
#1;data_in = testData6[2450];
@(posedge clk);
#1;data_in = testData6[2451];
@(posedge clk);
#1;data_in = testData6[2452];
@(posedge clk);
#1;data_in = testData6[2453];
@(posedge clk);
#1;data_in = testData6[2454];
@(posedge clk);
#1;data_in = testData6[2455];
@(posedge clk);
#1;data_in = testData6[2456];
@(posedge clk);
#1;data_in = testData6[2457];
@(posedge clk);
#1;data_in = testData6[2458];
@(posedge clk);
#1;data_in = testData6[2459];
@(posedge clk);
#1;data_in = testData6[2460];
@(posedge clk);
#1;data_in = testData6[2461];
@(posedge clk);
#1;data_in = testData6[2462];
@(posedge clk);
#1;data_in = testData6[2463];
@(posedge clk);
#1;data_in = testData6[2464];
@(posedge clk);
#1;data_in = testData6[2465];
@(posedge clk);
#1;data_in = testData6[2466];
@(posedge clk);
#1;data_in = testData6[2467];
@(posedge clk);
#1;data_in = testData6[2468];
@(posedge clk);
#1;data_in = testData6[2469];
@(posedge clk);
#1;data_in = testData6[2470];
@(posedge clk);
#1;data_in = testData6[2471];
@(posedge clk);
#1;data_in = testData6[2472];
@(posedge clk);
#1;data_in = testData6[2473];
@(posedge clk);
#1;data_in = testData6[2474];
@(posedge clk);
#1;data_in = testData6[2475];
@(posedge clk);
#1;data_in = testData6[2476];
@(posedge clk);
#1;data_in = testData6[2477];
@(posedge clk);
#1;data_in = testData6[2478];
@(posedge clk);
#1;data_in = testData6[2479];
@(posedge clk);
#1;data_in = testData6[2480];
@(posedge clk);
#1;data_in = testData6[2481];
@(posedge clk);
#1;data_in = testData6[2482];
@(posedge clk);
#1;data_in = testData6[2483];
@(posedge clk);
#1;data_in = testData6[2484];
@(posedge clk);
#1;data_in = testData6[2485];
@(posedge clk);
#1;data_in = testData6[2486];
@(posedge clk);
#1;data_in = testData6[2487];
@(posedge clk);
#1;data_in = testData6[2488];
@(posedge clk);
#1;data_in = testData6[2489];
@(posedge clk);
#1;data_in = testData6[2490];
@(posedge clk);
#1;data_in = testData6[2491];
@(posedge clk);
#1;data_in = testData6[2492];
@(posedge clk);
#1;data_in = testData6[2493];
@(posedge clk);
#1;data_in = testData6[2494];
@(posedge clk);
#1;data_in = testData6[2495];
@(posedge clk);
#1;data_in = testData6[2496];
@(posedge clk);
#1;data_in = testData6[2497];
@(posedge clk);
#1;data_in = testData6[2498];
@(posedge clk);
#1;data_in = testData6[2499];
@(posedge clk);
#1;data_in = testData6[2500];
@(posedge clk);
#1;data_in = testData6[2501];
@(posedge clk);
#1;data_in = testData6[2502];
@(posedge clk);
#1;data_in = testData6[2503];
@(posedge clk);
#1;data_in = testData6[2504];
@(posedge clk);
#1;data_in = testData6[2505];
@(posedge clk);
#1;data_in = testData6[2506];
@(posedge clk);
#1;data_in = testData6[2507];
@(posedge clk);
#1;data_in = testData6[2508];
@(posedge clk);
#1;data_in = testData6[2509];
@(posedge clk);
#1;data_in = testData6[2510];
@(posedge clk);
#1;data_in = testData6[2511];
@(posedge clk);
#1;data_in = testData6[2512];
@(posedge clk);
#1;data_in = testData6[2513];
@(posedge clk);
#1;data_in = testData6[2514];
@(posedge clk);
#1;data_in = testData6[2515];
@(posedge clk);
#1;data_in = testData6[2516];
@(posedge clk);
#1;data_in = testData6[2517];
@(posedge clk);
#1;data_in = testData6[2518];
@(posedge clk);
#1;data_in = testData6[2519];
@(posedge clk);
#1;data_in = testData6[2520];
@(posedge clk);
#1;data_in = testData6[2521];
@(posedge clk);
#1;data_in = testData6[2522];
@(posedge clk);
#1;data_in = testData6[2523];
@(posedge clk);
#1;data_in = testData6[2524];
@(posedge clk);
#1;data_in = testData6[2525];
@(posedge clk);
#1;data_in = testData6[2526];
@(posedge clk);
#1;data_in = testData6[2527];
@(posedge clk);
#1;data_in = testData6[2528];
@(posedge clk);
#1;data_in = testData6[2529];
@(posedge clk);
#1;data_in = testData6[2530];
@(posedge clk);
#1;data_in = testData6[2531];
@(posedge clk);
#1;data_in = testData6[2532];
@(posedge clk);
#1;data_in = testData6[2533];
@(posedge clk);
#1;data_in = testData6[2534];
@(posedge clk);
#1;data_in = testData6[2535];
@(posedge clk);
#1;data_in = testData6[2536];
@(posedge clk);
#1;data_in = testData6[2537];
@(posedge clk);
#1;data_in = testData6[2538];
@(posedge clk);
#1;data_in = testData6[2539];
@(posedge clk);
#1;data_in = testData6[2540];
@(posedge clk);
#1;data_in = testData6[2541];
@(posedge clk);
#1;data_in = testData6[2542];
@(posedge clk);
#1;data_in = testData6[2543];
@(posedge clk);
#1;data_in = testData6[2544];
@(posedge clk);
#1;data_in = testData6[2545];
@(posedge clk);
#1;data_in = testData6[2546];
@(posedge clk);
#1;data_in = testData6[2547];
@(posedge clk);
#1;data_in = testData6[2548];
@(posedge clk);
#1;data_in = testData6[2549];
@(posedge clk);
#1;data_in = testData6[2550];
@(posedge clk);
#1;data_in = testData6[2551];
@(posedge clk);
#1;data_in = testData6[2552];
@(posedge clk);
#1;data_in = testData6[2553];
@(posedge clk);
#1;data_in = testData6[2554];
@(posedge clk);
#1;data_in = testData6[2555];
@(posedge clk);
#1;data_in = testData6[2556];
@(posedge clk);
#1;data_in = testData6[2557];
@(posedge clk);
#1;data_in = testData6[2558];
@(posedge clk);
#1;data_in = testData6[2559];
@(posedge clk);
#1;data_in = testData6[2560];
@(posedge clk);
#1;data_in = testData6[2561];
@(posedge clk);
#1;data_in = testData6[2562];
@(posedge clk);
#1;data_in = testData6[2563];
@(posedge clk);
#1;data_in = testData6[2564];
@(posedge clk);
#1;data_in = testData6[2565];
@(posedge clk);
#1;data_in = testData6[2566];
@(posedge clk);
#1;data_in = testData6[2567];
@(posedge clk);
#1;data_in = testData6[2568];
@(posedge clk);
#1;data_in = testData6[2569];
@(posedge clk);
#1;data_in = testData6[2570];
@(posedge clk);
#1;data_in = testData6[2571];
@(posedge clk);
#1;data_in = testData6[2572];
@(posedge clk);
#1;data_in = testData6[2573];
@(posedge clk);
#1;data_in = testData6[2574];
@(posedge clk);
#1;data_in = testData6[2575];
@(posedge clk);
#1;data_in = testData6[2576];
@(posedge clk);
#1;data_in = testData6[2577];
@(posedge clk);
#1;data_in = testData6[2578];
@(posedge clk);
#1;data_in = testData6[2579];
@(posedge clk);
#1;data_in = testData6[2580];
@(posedge clk);
#1;data_in = testData6[2581];
@(posedge clk);
#1;data_in = testData6[2582];
@(posedge clk);
#1;data_in = testData6[2583];
@(posedge clk);
#1;data_in = testData6[2584];
@(posedge clk);
#1;data_in = testData6[2585];
@(posedge clk);
#1;data_in = testData6[2586];
@(posedge clk);
#1;data_in = testData6[2587];
@(posedge clk);
#1;data_in = testData6[2588];
@(posedge clk);
#1;data_in = testData6[2589];
@(posedge clk);
#1;data_in = testData6[2590];
@(posedge clk);
#1;data_in = testData6[2591];
@(posedge clk);
#1;data_in = testData6[2592];
@(posedge clk);
#1;data_in = testData6[2593];
@(posedge clk);
#1;data_in = testData6[2594];
@(posedge clk);
#1;data_in = testData6[2595];
@(posedge clk);
#1;data_in = testData6[2596];
@(posedge clk);
#1;data_in = testData6[2597];
@(posedge clk);
#1;data_in = testData6[2598];
@(posedge clk);
#1;data_in = testData6[2599];
@(posedge clk);
#1;data_in = testData6[2600];
@(posedge clk);
#1;data_in = testData6[2601];
@(posedge clk);
#1;data_in = testData6[2602];
@(posedge clk);
#1;data_in = testData6[2603];
@(posedge clk);
#1;data_in = testData6[2604];
@(posedge clk);
#1;data_in = testData6[2605];
@(posedge clk);
#1;data_in = testData6[2606];
@(posedge clk);
#1;data_in = testData6[2607];
@(posedge clk);
#1;data_in = testData6[2608];
@(posedge clk);
#1;data_in = testData6[2609];
@(posedge clk);
#1;data_in = testData6[2610];
@(posedge clk);
#1;data_in = testData6[2611];
@(posedge clk);
#1;data_in = testData6[2612];
@(posedge clk);
#1;data_in = testData6[2613];
@(posedge clk);
#1;data_in = testData6[2614];
@(posedge clk);
#1;data_in = testData6[2615];
@(posedge clk);
#1;data_in = testData6[2616];
@(posedge clk);
#1;data_in = testData6[2617];
@(posedge clk);
#1;data_in = testData6[2618];
@(posedge clk);
#1;data_in = testData6[2619];
@(posedge clk);
#1;data_in = testData6[2620];
@(posedge clk);
#1;data_in = testData6[2621];
@(posedge clk);
#1;data_in = testData6[2622];
@(posedge clk);
#1;data_in = testData6[2623];
@(posedge clk);
#1;data_in = testData6[2624];
@(posedge clk);
#1;data_in = testData6[2625];
@(posedge clk);
#1;data_in = testData6[2626];
@(posedge clk);
#1;data_in = testData6[2627];
@(posedge clk);
#1;data_in = testData6[2628];
@(posedge clk);
#1;data_in = testData6[2629];
@(posedge clk);
#1;data_in = testData6[2630];
@(posedge clk);
#1;data_in = testData6[2631];
@(posedge clk);
#1;data_in = testData6[2632];
@(posedge clk);
#1;data_in = testData6[2633];
@(posedge clk);
#1;data_in = testData6[2634];
@(posedge clk);
#1;data_in = testData6[2635];
@(posedge clk);
#1;data_in = testData6[2636];
@(posedge clk);
#1;data_in = testData6[2637];
@(posedge clk);
#1;data_in = testData6[2638];
@(posedge clk);
#1;data_in = testData6[2639];
@(posedge clk);
#1;data_in = testData6[2640];
@(posedge clk);
#1;data_in = testData6[2641];
@(posedge clk);
#1;data_in = testData6[2642];
@(posedge clk);
#1;data_in = testData6[2643];
@(posedge clk);
#1;data_in = testData6[2644];
@(posedge clk);
#1;data_in = testData6[2645];
@(posedge clk);
#1;data_in = testData6[2646];
@(posedge clk);
#1;data_in = testData6[2647];
@(posedge clk);
#1;data_in = testData6[2648];
@(posedge clk);
#1;data_in = testData6[2649];
@(posedge clk);
#1;data_in = testData6[2650];
@(posedge clk);
#1;data_in = testData6[2651];
@(posedge clk);
#1;data_in = testData6[2652];
@(posedge clk);
#1;data_in = testData6[2653];
@(posedge clk);
#1;data_in = testData6[2654];
@(posedge clk);
#1;data_in = testData6[2655];
@(posedge clk);
#1;data_in = testData6[2656];
@(posedge clk);
#1;data_in = testData6[2657];
@(posedge clk);
#1;data_in = testData6[2658];
@(posedge clk);
#1;data_in = testData6[2659];
@(posedge clk);
#1;data_in = testData6[2660];
@(posedge clk);
#1;data_in = testData6[2661];
@(posedge clk);
#1;data_in = testData6[2662];
@(posedge clk);
#1;data_in = testData6[2663];
@(posedge clk);
#1;data_in = testData6[2664];
@(posedge clk);
#1;data_in = testData6[2665];
@(posedge clk);
#1;data_in = testData6[2666];
@(posedge clk);
#1;data_in = testData6[2667];
@(posedge clk);
#1;data_in = testData6[2668];
@(posedge clk);
#1;data_in = testData6[2669];
@(posedge clk);
#1;data_in = testData6[2670];
@(posedge clk);
#1;data_in = testData6[2671];
@(posedge clk);
#1;data_in = testData6[2672];
@(posedge clk);
#1;data_in = testData6[2673];
@(posedge clk);
#1;data_in = testData6[2674];
@(posedge clk);
#1;data_in = testData6[2675];
@(posedge clk);
#1;data_in = testData6[2676];
@(posedge clk);
#1;data_in = testData6[2677];
@(posedge clk);
#1;data_in = testData6[2678];
@(posedge clk);
#1;data_in = testData6[2679];
@(posedge clk);
#1;data_in = testData6[2680];
@(posedge clk);
#1;data_in = testData6[2681];
@(posedge clk);
#1;data_in = testData6[2682];
@(posedge clk);
#1;data_in = testData6[2683];
@(posedge clk);
#1;data_in = testData6[2684];
@(posedge clk);
#1;data_in = testData6[2685];
@(posedge clk);
#1;data_in = testData6[2686];
@(posedge clk);
#1;data_in = testData6[2687];
@(posedge clk);
#1;data_in = testData6[2688];
@(posedge clk);
#1;data_in = testData6[2689];
@(posedge clk);
#1;data_in = testData6[2690];
@(posedge clk);
#1;data_in = testData6[2691];
@(posedge clk);
#1;data_in = testData6[2692];
@(posedge clk);
#1;data_in = testData6[2693];
@(posedge clk);
#1;data_in = testData6[2694];
@(posedge clk);
#1;data_in = testData6[2695];
@(posedge clk);
#1;data_in = testData6[2696];
@(posedge clk);
#1;data_in = testData6[2697];
@(posedge clk);
#1;data_in = testData6[2698];
@(posedge clk);
#1;data_in = testData6[2699];
@(posedge clk);
#1;data_in = testData6[2700];
@(posedge clk);
#1;data_in = testData6[2701];
@(posedge clk);
#1;data_in = testData6[2702];
@(posedge clk);
#1;data_in = testData6[2703];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2704]; 
@(posedge clk);
#1;data_in = testData6[2705];
@(posedge clk);
#1;data_in = testData6[2706];
@(posedge clk);
#1;data_in = testData6[2707];
@(posedge clk);
#1;data_in = testData6[2708];
@(posedge clk);
#1;data_in = testData6[2709];
@(posedge clk);
#1;data_in = testData6[2710];
@(posedge clk);
#1;data_in = testData6[2711];
@(posedge clk);
#1;data_in = testData6[2712];
@(posedge clk);
#1;data_in = testData6[2713];
@(posedge clk);
#1;data_in = testData6[2714];
@(posedge clk);
#1;data_in = testData6[2715];
@(posedge clk);
#1;data_in = testData6[2716];
@(posedge clk);
#1;data_in = testData6[2717];
@(posedge clk);
#1;data_in = testData6[2718];
@(posedge clk);
#1;data_in = testData6[2719];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2720];
@(posedge clk);
#1;data_in = testData6[2721];
@(posedge clk);
#1;data_in = testData6[2722];
@(posedge clk);
#1;data_in = testData6[2723];
@(posedge clk);
#1;data_in = testData6[2724];
@(posedge clk);
#1;data_in = testData6[2725];
@(posedge clk);
#1;data_in = testData6[2726];
@(posedge clk);
#1;data_in = testData6[2727];
@(posedge clk);
#1;data_in = testData6[2728];
@(posedge clk);
#1;data_in = testData6[2729];
@(posedge clk);
#1;data_in = testData6[2730];
@(posedge clk);
#1;data_in = testData6[2731];
@(posedge clk);
#1;data_in = testData6[2732];
@(posedge clk);
#1;data_in = testData6[2733];
@(posedge clk);
#1;data_in = testData6[2734];
@(posedge clk);
#1;data_in = testData6[2735];
@(posedge clk);
#1;data_in = testData6[2736];
@(posedge clk);
#1;data_in = testData6[2737];
@(posedge clk);
#1;data_in = testData6[2738];
@(posedge clk);
#1;data_in = testData6[2739];
@(posedge clk);
#1;data_in = testData6[2740];
@(posedge clk);
#1;data_in = testData6[2741];
@(posedge clk);
#1;data_in = testData6[2742];
@(posedge clk);
#1;data_in = testData6[2743];
@(posedge clk);
#1;data_in = testData6[2744];
@(posedge clk);
#1;data_in = testData6[2745];
@(posedge clk);
#1;data_in = testData6[2746];
@(posedge clk);
#1;data_in = testData6[2747];
@(posedge clk);
#1;data_in = testData6[2748];
@(posedge clk);
#1;data_in = testData6[2749];
@(posedge clk);
#1;data_in = testData6[2750];
@(posedge clk);
#1;data_in = testData6[2751];
@(posedge clk);
#1;data_in = testData6[2752];
@(posedge clk);
#1;data_in = testData6[2753];
@(posedge clk);
#1;data_in = testData6[2754];
@(posedge clk);
#1;data_in = testData6[2755];
@(posedge clk);
#1;data_in = testData6[2756];
@(posedge clk);
#1;data_in = testData6[2757];
@(posedge clk);
#1;data_in = testData6[2758];
@(posedge clk);
#1;data_in = testData6[2759];
@(posedge clk);
#1;data_in = testData6[2760];
@(posedge clk);
#1;data_in = testData6[2761];
@(posedge clk);
#1;data_in = testData6[2762];
@(posedge clk);
#1;data_in = testData6[2763];
@(posedge clk);
#1;data_in = testData6[2764];
@(posedge clk);
#1;data_in = testData6[2765];
@(posedge clk);
#1;data_in = testData6[2766];
@(posedge clk);
#1;data_in = testData6[2767];
@(posedge clk);
#1;data_in = testData6[2768];
@(posedge clk);
#1;data_in = testData6[2769];
@(posedge clk);
#1;data_in = testData6[2770];
@(posedge clk);
#1;data_in = testData6[2771];
@(posedge clk);
#1;data_in = testData6[2772];
@(posedge clk);
#1;data_in = testData6[2773];
@(posedge clk);
#1;data_in = testData6[2774];
@(posedge clk);
#1;data_in = testData6[2775];
@(posedge clk);
#1;data_in = testData6[2776];
@(posedge clk);
#1;data_in = testData6[2777];
@(posedge clk);
#1;data_in = testData6[2778];
@(posedge clk);
#1;data_in = testData6[2779];
@(posedge clk);
#1;data_in = testData6[2780];
@(posedge clk);
#1;data_in = testData6[2781];
@(posedge clk);
#1;data_in = testData6[2782];
@(posedge clk);
#1;data_in = testData6[2783];
@(posedge clk);
#1;data_in = testData6[2784];
@(posedge clk);
#1;data_in = testData6[2785];
@(posedge clk);
#1;data_in = testData6[2786];
@(posedge clk);
#1;data_in = testData6[2787];
@(posedge clk);
#1;data_in = testData6[2788];
@(posedge clk);
#1;data_in = testData6[2789];
@(posedge clk);
#1;data_in = testData6[2790];
@(posedge clk);
#1;data_in = testData6[2791];
@(posedge clk);
#1;data_in = testData6[2792];
@(posedge clk);
#1;data_in = testData6[2793];
@(posedge clk);
#1;data_in = testData6[2794];
@(posedge clk);
#1;data_in = testData6[2795];
@(posedge clk);
#1;data_in = testData6[2796];
@(posedge clk);
#1;data_in = testData6[2797];
@(posedge clk);
#1;data_in = testData6[2798];
@(posedge clk);
#1;data_in = testData6[2799];
@(posedge clk);
#1;data_in = testData6[2800];
@(posedge clk);
#1;data_in = testData6[2801];
@(posedge clk);
#1;data_in = testData6[2802];
@(posedge clk);
#1;data_in = testData6[2803];
@(posedge clk);
#1;data_in = testData6[2804];
@(posedge clk);
#1;data_in = testData6[2805];
@(posedge clk);
#1;data_in = testData6[2806];
@(posedge clk);
#1;data_in = testData6[2807];
@(posedge clk);
#1;data_in = testData6[2808];
@(posedge clk);
#1;data_in = testData6[2809];
@(posedge clk);
#1;data_in = testData6[2810];
@(posedge clk);
#1;data_in = testData6[2811];
@(posedge clk);
#1;data_in = testData6[2812];
@(posedge clk);
#1;data_in = testData6[2813];
@(posedge clk);
#1;data_in = testData6[2814];
@(posedge clk);
#1;data_in = testData6[2815];
@(posedge clk);
#1;data_in = testData6[2816];
@(posedge clk);
#1;data_in = testData6[2817];
@(posedge clk);
#1;data_in = testData6[2818];
@(posedge clk);
#1;data_in = testData6[2819];
@(posedge clk);
#1;data_in = testData6[2820];
@(posedge clk);
#1;data_in = testData6[2821];
@(posedge clk);
#1;data_in = testData6[2822];
@(posedge clk);
#1;data_in = testData6[2823];
@(posedge clk);
#1;data_in = testData6[2824];
@(posedge clk);
#1;data_in = testData6[2825];
@(posedge clk);
#1;data_in = testData6[2826];
@(posedge clk);
#1;data_in = testData6[2827];
@(posedge clk);
#1;data_in = testData6[2828];
@(posedge clk);
#1;data_in = testData6[2829];
@(posedge clk);
#1;data_in = testData6[2830];
@(posedge clk);
#1;data_in = testData6[2831];
@(posedge clk);
#1;data_in = testData6[2832];
@(posedge clk);
#1;data_in = testData6[2833];
@(posedge clk);
#1;data_in = testData6[2834];
@(posedge clk);
#1;data_in = testData6[2835];
@(posedge clk);
#1;data_in = testData6[2836];
@(posedge clk);
#1;data_in = testData6[2837];
@(posedge clk);
#1;data_in = testData6[2838];
@(posedge clk);
#1;data_in = testData6[2839];
@(posedge clk);
#1;data_in = testData6[2840];
@(posedge clk);
#1;data_in = testData6[2841];
@(posedge clk);
#1;data_in = testData6[2842];
@(posedge clk);
#1;data_in = testData6[2843];
@(posedge clk);
#1;data_in = testData6[2844];
@(posedge clk);
#1;data_in = testData6[2845];
@(posedge clk);
#1;data_in = testData6[2846];
@(posedge clk);
#1;data_in = testData6[2847];
@(posedge clk);
#1;data_in = testData6[2848];
@(posedge clk);
#1;data_in = testData6[2849];
@(posedge clk);
#1;data_in = testData6[2850];
@(posedge clk);
#1;data_in = testData6[2851];
@(posedge clk);
#1;data_in = testData6[2852];
@(posedge clk);
#1;data_in = testData6[2853];
@(posedge clk);
#1;data_in = testData6[2854];
@(posedge clk);
#1;data_in = testData6[2855];
@(posedge clk);
#1;data_in = testData6[2856];
@(posedge clk);
#1;data_in = testData6[2857];
@(posedge clk);
#1;data_in = testData6[2858];
@(posedge clk);
#1;data_in = testData6[2859];
@(posedge clk);
#1;data_in = testData6[2860];
@(posedge clk);
#1;data_in = testData6[2861];
@(posedge clk);
#1;data_in = testData6[2862];
@(posedge clk);
#1;data_in = testData6[2863];
@(posedge clk);
#1;data_in = testData6[2864];
@(posedge clk);
#1;data_in = testData6[2865];
@(posedge clk);
#1;data_in = testData6[2866];
@(posedge clk);
#1;data_in = testData6[2867];
@(posedge clk);
#1;data_in = testData6[2868];
@(posedge clk);
#1;data_in = testData6[2869];
@(posedge clk);
#1;data_in = testData6[2870];
@(posedge clk);
#1;data_in = testData6[2871];
@(posedge clk);
#1;data_in = testData6[2872];
@(posedge clk);
#1;data_in = testData6[2873];
@(posedge clk);
#1;data_in = testData6[2874];
@(posedge clk);
#1;data_in = testData6[2875];
@(posedge clk);
#1;data_in = testData6[2876];
@(posedge clk);
#1;data_in = testData6[2877];
@(posedge clk);
#1;data_in = testData6[2878];
@(posedge clk);
#1;data_in = testData6[2879];
@(posedge clk);
#1;data_in = testData6[2880];
@(posedge clk);
#1;data_in = testData6[2881];
@(posedge clk);
#1;data_in = testData6[2882];
@(posedge clk);
#1;data_in = testData6[2883];
@(posedge clk);
#1;data_in = testData6[2884];
@(posedge clk);
#1;data_in = testData6[2885];
@(posedge clk);
#1;data_in = testData6[2886];
@(posedge clk);
#1;data_in = testData6[2887];
@(posedge clk);
#1;data_in = testData6[2888];
@(posedge clk);
#1;data_in = testData6[2889];
@(posedge clk);
#1;data_in = testData6[2890];
@(posedge clk);
#1;data_in = testData6[2891];
@(posedge clk);
#1;data_in = testData6[2892];
@(posedge clk);
#1;data_in = testData6[2893];
@(posedge clk);
#1;data_in = testData6[2894];
@(posedge clk);
#1;data_in = testData6[2895];
@(posedge clk);
#1;data_in = testData6[2896];
@(posedge clk);
#1;data_in = testData6[2897];
@(posedge clk);
#1;data_in = testData6[2898];
@(posedge clk);
#1;data_in = testData6[2899];
@(posedge clk);
#1;data_in = testData6[2900];
@(posedge clk);
#1;data_in = testData6[2901];
@(posedge clk);
#1;data_in = testData6[2902];
@(posedge clk);
#1;data_in = testData6[2903];
@(posedge clk);
#1;data_in = testData6[2904];
@(posedge clk);
#1;data_in = testData6[2905];
@(posedge clk);
#1;data_in = testData6[2906];
@(posedge clk);
#1;data_in = testData6[2907];
@(posedge clk);
#1;data_in = testData6[2908];
@(posedge clk);
#1;data_in = testData6[2909];
@(posedge clk);
#1;data_in = testData6[2910];
@(posedge clk);
#1;data_in = testData6[2911];
@(posedge clk);
#1;data_in = testData6[2912];
@(posedge clk);
#1;data_in = testData6[2913];
@(posedge clk);
#1;data_in = testData6[2914];
@(posedge clk);
#1;data_in = testData6[2915];
@(posedge clk);
#1;data_in = testData6[2916];
@(posedge clk);
#1;data_in = testData6[2917];
@(posedge clk);
#1;data_in = testData6[2918];
@(posedge clk);
#1;data_in = testData6[2919];
@(posedge clk);
#1;data_in = testData6[2920];
@(posedge clk);
#1;data_in = testData6[2921];
@(posedge clk);
#1;data_in = testData6[2922];
@(posedge clk);
#1;data_in = testData6[2923];
@(posedge clk);
#1;data_in = testData6[2924];
@(posedge clk);
#1;data_in = testData6[2925];
@(posedge clk);
#1;data_in = testData6[2926];
@(posedge clk);
#1;data_in = testData6[2927];
@(posedge clk);
#1;data_in = testData6[2928];
@(posedge clk);
#1;data_in = testData6[2929];
@(posedge clk);
#1;data_in = testData6[2930];
@(posedge clk);
#1;data_in = testData6[2931];
@(posedge clk);
#1;data_in = testData6[2932];
@(posedge clk);
#1;data_in = testData6[2933];
@(posedge clk);
#1;data_in = testData6[2934];
@(posedge clk);
#1;data_in = testData6[2935];
@(posedge clk);
#1;data_in = testData6[2936];
@(posedge clk);
#1;data_in = testData6[2937];
@(posedge clk);
#1;data_in = testData6[2938];
@(posedge clk);
#1;data_in = testData6[2939];
@(posedge clk);
#1;data_in = testData6[2940];
@(posedge clk);
#1;data_in = testData6[2941];
@(posedge clk);
#1;data_in = testData6[2942];
@(posedge clk);
#1;data_in = testData6[2943];
@(posedge clk);
#1;data_in = testData6[2944];
@(posedge clk);
#1;data_in = testData6[2945];
@(posedge clk);
#1;data_in = testData6[2946];
@(posedge clk);
#1;data_in = testData6[2947];
@(posedge clk);
#1;data_in = testData6[2948];
@(posedge clk);
#1;data_in = testData6[2949];
@(posedge clk);
#1;data_in = testData6[2950];
@(posedge clk);
#1;data_in = testData6[2951];
@(posedge clk);
#1;data_in = testData6[2952];
@(posedge clk);
#1;data_in = testData6[2953];
@(posedge clk);
#1;data_in = testData6[2954];
@(posedge clk);
#1;data_in = testData6[2955];
@(posedge clk);
#1;data_in = testData6[2956];
@(posedge clk);
#1;data_in = testData6[2957];
@(posedge clk);
#1;data_in = testData6[2958];
@(posedge clk);
#1;data_in = testData6[2959];
@(posedge clk);
#1;data_in = testData6[2960];
@(posedge clk);
#1;data_in = testData6[2961];
@(posedge clk);
#1;data_in = testData6[2962];
@(posedge clk);
#1;data_in = testData6[2963];
@(posedge clk);
#1;data_in = testData6[2964];
@(posedge clk);
#1;data_in = testData6[2965];
@(posedge clk);
#1;data_in = testData6[2966];
@(posedge clk);
#1;data_in = testData6[2967];
@(posedge clk);
#1;data_in = testData6[2968];
@(posedge clk);
#1;data_in = testData6[2969];
@(posedge clk);
#1;data_in = testData6[2970];
@(posedge clk);
#1;data_in = testData6[2971];
@(posedge clk);
#1;data_in = testData6[2972];
@(posedge clk);
#1;data_in = testData6[2973];
@(posedge clk);
#1;data_in = testData6[2974];
@(posedge clk);
#1;data_in = testData6[2975];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2976]; 
@(posedge clk);
#1;data_in = testData6[2977];
@(posedge clk);
#1;data_in = testData6[2978];
@(posedge clk);
#1;data_in = testData6[2979];
@(posedge clk);
#1;data_in = testData6[2980];
@(posedge clk);
#1;data_in = testData6[2981];
@(posedge clk);
#1;data_in = testData6[2982];
@(posedge clk);
#1;data_in = testData6[2983];
@(posedge clk);
#1;data_in = testData6[2984];
@(posedge clk);
#1;data_in = testData6[2985];
@(posedge clk);
#1;data_in = testData6[2986];
@(posedge clk);
#1;data_in = testData6[2987];
@(posedge clk);
#1;data_in = testData6[2988];
@(posedge clk);
#1;data_in = testData6[2989];
@(posedge clk);
#1;data_in = testData6[2990];
@(posedge clk);
#1;data_in = testData6[2991];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2992];
@(posedge clk);
#1;data_in = testData6[2993];
@(posedge clk);
#1;data_in = testData6[2994];
@(posedge clk);
#1;data_in = testData6[2995];
@(posedge clk);
#1;data_in = testData6[2996];
@(posedge clk);
#1;data_in = testData6[2997];
@(posedge clk);
#1;data_in = testData6[2998];
@(posedge clk);
#1;data_in = testData6[2999];
@(posedge clk);
#1;data_in = testData6[3000];
@(posedge clk);
#1;data_in = testData6[3001];
@(posedge clk);
#1;data_in = testData6[3002];
@(posedge clk);
#1;data_in = testData6[3003];
@(posedge clk);
#1;data_in = testData6[3004];
@(posedge clk);
#1;data_in = testData6[3005];
@(posedge clk);
#1;data_in = testData6[3006];
@(posedge clk);
#1;data_in = testData6[3007];
@(posedge clk);
#1;data_in = testData6[3008];
@(posedge clk);
#1;data_in = testData6[3009];
@(posedge clk);
#1;data_in = testData6[3010];
@(posedge clk);
#1;data_in = testData6[3011];
@(posedge clk);
#1;data_in = testData6[3012];
@(posedge clk);
#1;data_in = testData6[3013];
@(posedge clk);
#1;data_in = testData6[3014];
@(posedge clk);
#1;data_in = testData6[3015];
@(posedge clk);
#1;data_in = testData6[3016];
@(posedge clk);
#1;data_in = testData6[3017];
@(posedge clk);
#1;data_in = testData6[3018];
@(posedge clk);
#1;data_in = testData6[3019];
@(posedge clk);
#1;data_in = testData6[3020];
@(posedge clk);
#1;data_in = testData6[3021];
@(posedge clk);
#1;data_in = testData6[3022];
@(posedge clk);
#1;data_in = testData6[3023];
@(posedge clk);
#1;data_in = testData6[3024];
@(posedge clk);
#1;data_in = testData6[3025];
@(posedge clk);
#1;data_in = testData6[3026];
@(posedge clk);
#1;data_in = testData6[3027];
@(posedge clk);
#1;data_in = testData6[3028];
@(posedge clk);
#1;data_in = testData6[3029];
@(posedge clk);
#1;data_in = testData6[3030];
@(posedge clk);
#1;data_in = testData6[3031];
@(posedge clk);
#1;data_in = testData6[3032];
@(posedge clk);
#1;data_in = testData6[3033];
@(posedge clk);
#1;data_in = testData6[3034];
@(posedge clk);
#1;data_in = testData6[3035];
@(posedge clk);
#1;data_in = testData6[3036];
@(posedge clk);
#1;data_in = testData6[3037];
@(posedge clk);
#1;data_in = testData6[3038];
@(posedge clk);
#1;data_in = testData6[3039];
@(posedge clk);
#1;data_in = testData6[3040];
@(posedge clk);
#1;data_in = testData6[3041];
@(posedge clk);
#1;data_in = testData6[3042];
@(posedge clk);
#1;data_in = testData6[3043];
@(posedge clk);
#1;data_in = testData6[3044];
@(posedge clk);
#1;data_in = testData6[3045];
@(posedge clk);
#1;data_in = testData6[3046];
@(posedge clk);
#1;data_in = testData6[3047];
@(posedge clk);
#1;data_in = testData6[3048];
@(posedge clk);
#1;data_in = testData6[3049];
@(posedge clk);
#1;data_in = testData6[3050];
@(posedge clk);
#1;data_in = testData6[3051];
@(posedge clk);
#1;data_in = testData6[3052];
@(posedge clk);
#1;data_in = testData6[3053];
@(posedge clk);
#1;data_in = testData6[3054];
@(posedge clk);
#1;data_in = testData6[3055];
@(posedge clk);
#1;data_in = testData6[3056];
@(posedge clk);
#1;data_in = testData6[3057];
@(posedge clk);
#1;data_in = testData6[3058];
@(posedge clk);
#1;data_in = testData6[3059];
@(posedge clk);
#1;data_in = testData6[3060];
@(posedge clk);
#1;data_in = testData6[3061];
@(posedge clk);
#1;data_in = testData6[3062];
@(posedge clk);
#1;data_in = testData6[3063];
@(posedge clk);
#1;data_in = testData6[3064];
@(posedge clk);
#1;data_in = testData6[3065];
@(posedge clk);
#1;data_in = testData6[3066];
@(posedge clk);
#1;data_in = testData6[3067];
@(posedge clk);
#1;data_in = testData6[3068];
@(posedge clk);
#1;data_in = testData6[3069];
@(posedge clk);
#1;data_in = testData6[3070];
@(posedge clk);
#1;data_in = testData6[3071];
@(posedge clk);
#1;data_in = testData6[3072];
@(posedge clk);
#1;data_in = testData6[3073];
@(posedge clk);
#1;data_in = testData6[3074];
@(posedge clk);
#1;data_in = testData6[3075];
@(posedge clk);
#1;data_in = testData6[3076];
@(posedge clk);
#1;data_in = testData6[3077];
@(posedge clk);
#1;data_in = testData6[3078];
@(posedge clk);
#1;data_in = testData6[3079];
@(posedge clk);
#1;data_in = testData6[3080];
@(posedge clk);
#1;data_in = testData6[3081];
@(posedge clk);
#1;data_in = testData6[3082];
@(posedge clk);
#1;data_in = testData6[3083];
@(posedge clk);
#1;data_in = testData6[3084];
@(posedge clk);
#1;data_in = testData6[3085];
@(posedge clk);
#1;data_in = testData6[3086];
@(posedge clk);
#1;data_in = testData6[3087];
@(posedge clk);
#1;data_in = testData6[3088];
@(posedge clk);
#1;data_in = testData6[3089];
@(posedge clk);
#1;data_in = testData6[3090];
@(posedge clk);
#1;data_in = testData6[3091];
@(posedge clk);
#1;data_in = testData6[3092];
@(posedge clk);
#1;data_in = testData6[3093];
@(posedge clk);
#1;data_in = testData6[3094];
@(posedge clk);
#1;data_in = testData6[3095];
@(posedge clk);
#1;data_in = testData6[3096];
@(posedge clk);
#1;data_in = testData6[3097];
@(posedge clk);
#1;data_in = testData6[3098];
@(posedge clk);
#1;data_in = testData6[3099];
@(posedge clk);
#1;data_in = testData6[3100];
@(posedge clk);
#1;data_in = testData6[3101];
@(posedge clk);
#1;data_in = testData6[3102];
@(posedge clk);
#1;data_in = testData6[3103];
@(posedge clk);
#1;data_in = testData6[3104];
@(posedge clk);
#1;data_in = testData6[3105];
@(posedge clk);
#1;data_in = testData6[3106];
@(posedge clk);
#1;data_in = testData6[3107];
@(posedge clk);
#1;data_in = testData6[3108];
@(posedge clk);
#1;data_in = testData6[3109];
@(posedge clk);
#1;data_in = testData6[3110];
@(posedge clk);
#1;data_in = testData6[3111];
@(posedge clk);
#1;data_in = testData6[3112];
@(posedge clk);
#1;data_in = testData6[3113];
@(posedge clk);
#1;data_in = testData6[3114];
@(posedge clk);
#1;data_in = testData6[3115];
@(posedge clk);
#1;data_in = testData6[3116];
@(posedge clk);
#1;data_in = testData6[3117];
@(posedge clk);
#1;data_in = testData6[3118];
@(posedge clk);
#1;data_in = testData6[3119];
@(posedge clk);
#1;data_in = testData6[3120];
@(posedge clk);
#1;data_in = testData6[3121];
@(posedge clk);
#1;data_in = testData6[3122];
@(posedge clk);
#1;data_in = testData6[3123];
@(posedge clk);
#1;data_in = testData6[3124];
@(posedge clk);
#1;data_in = testData6[3125];
@(posedge clk);
#1;data_in = testData6[3126];
@(posedge clk);
#1;data_in = testData6[3127];
@(posedge clk);
#1;data_in = testData6[3128];
@(posedge clk);
#1;data_in = testData6[3129];
@(posedge clk);
#1;data_in = testData6[3130];
@(posedge clk);
#1;data_in = testData6[3131];
@(posedge clk);
#1;data_in = testData6[3132];
@(posedge clk);
#1;data_in = testData6[3133];
@(posedge clk);
#1;data_in = testData6[3134];
@(posedge clk);
#1;data_in = testData6[3135];
@(posedge clk);
#1;data_in = testData6[3136];
@(posedge clk);
#1;data_in = testData6[3137];
@(posedge clk);
#1;data_in = testData6[3138];
@(posedge clk);
#1;data_in = testData6[3139];
@(posedge clk);
#1;data_in = testData6[3140];
@(posedge clk);
#1;data_in = testData6[3141];
@(posedge clk);
#1;data_in = testData6[3142];
@(posedge clk);
#1;data_in = testData6[3143];
@(posedge clk);
#1;data_in = testData6[3144];
@(posedge clk);
#1;data_in = testData6[3145];
@(posedge clk);
#1;data_in = testData6[3146];
@(posedge clk);
#1;data_in = testData6[3147];
@(posedge clk);
#1;data_in = testData6[3148];
@(posedge clk);
#1;data_in = testData6[3149];
@(posedge clk);
#1;data_in = testData6[3150];
@(posedge clk);
#1;data_in = testData6[3151];
@(posedge clk);
#1;data_in = testData6[3152];
@(posedge clk);
#1;data_in = testData6[3153];
@(posedge clk);
#1;data_in = testData6[3154];
@(posedge clk);
#1;data_in = testData6[3155];
@(posedge clk);
#1;data_in = testData6[3156];
@(posedge clk);
#1;data_in = testData6[3157];
@(posedge clk);
#1;data_in = testData6[3158];
@(posedge clk);
#1;data_in = testData6[3159];
@(posedge clk);
#1;data_in = testData6[3160];
@(posedge clk);
#1;data_in = testData6[3161];
@(posedge clk);
#1;data_in = testData6[3162];
@(posedge clk);
#1;data_in = testData6[3163];
@(posedge clk);
#1;data_in = testData6[3164];
@(posedge clk);
#1;data_in = testData6[3165];
@(posedge clk);
#1;data_in = testData6[3166];
@(posedge clk);
#1;data_in = testData6[3167];
@(posedge clk);
#1;data_in = testData6[3168];
@(posedge clk);
#1;data_in = testData6[3169];
@(posedge clk);
#1;data_in = testData6[3170];
@(posedge clk);
#1;data_in = testData6[3171];
@(posedge clk);
#1;data_in = testData6[3172];
@(posedge clk);
#1;data_in = testData6[3173];
@(posedge clk);
#1;data_in = testData6[3174];
@(posedge clk);
#1;data_in = testData6[3175];
@(posedge clk);
#1;data_in = testData6[3176];
@(posedge clk);
#1;data_in = testData6[3177];
@(posedge clk);
#1;data_in = testData6[3178];
@(posedge clk);
#1;data_in = testData6[3179];
@(posedge clk);
#1;data_in = testData6[3180];
@(posedge clk);
#1;data_in = testData6[3181];
@(posedge clk);
#1;data_in = testData6[3182];
@(posedge clk);
#1;data_in = testData6[3183];
@(posedge clk);
#1;data_in = testData6[3184];
@(posedge clk);
#1;data_in = testData6[3185];
@(posedge clk);
#1;data_in = testData6[3186];
@(posedge clk);
#1;data_in = testData6[3187];
@(posedge clk);
#1;data_in = testData6[3188];
@(posedge clk);
#1;data_in = testData6[3189];
@(posedge clk);
#1;data_in = testData6[3190];
@(posedge clk);
#1;data_in = testData6[3191];
@(posedge clk);
#1;data_in = testData6[3192];
@(posedge clk);
#1;data_in = testData6[3193];
@(posedge clk);
#1;data_in = testData6[3194];
@(posedge clk);
#1;data_in = testData6[3195];
@(posedge clk);
#1;data_in = testData6[3196];
@(posedge clk);
#1;data_in = testData6[3197];
@(posedge clk);
#1;data_in = testData6[3198];
@(posedge clk);
#1;data_in = testData6[3199];
@(posedge clk);
#1;data_in = testData6[3200];
@(posedge clk);
#1;data_in = testData6[3201];
@(posedge clk);
#1;data_in = testData6[3202];
@(posedge clk);
#1;data_in = testData6[3203];
@(posedge clk);
#1;data_in = testData6[3204];
@(posedge clk);
#1;data_in = testData6[3205];
@(posedge clk);
#1;data_in = testData6[3206];
@(posedge clk);
#1;data_in = testData6[3207];
@(posedge clk);
#1;data_in = testData6[3208];
@(posedge clk);
#1;data_in = testData6[3209];
@(posedge clk);
#1;data_in = testData6[3210];
@(posedge clk);
#1;data_in = testData6[3211];
@(posedge clk);
#1;data_in = testData6[3212];
@(posedge clk);
#1;data_in = testData6[3213];
@(posedge clk);
#1;data_in = testData6[3214];
@(posedge clk);
#1;data_in = testData6[3215];
@(posedge clk);
#1;data_in = testData6[3216];
@(posedge clk);
#1;data_in = testData6[3217];
@(posedge clk);
#1;data_in = testData6[3218];
@(posedge clk);
#1;data_in = testData6[3219];
@(posedge clk);
#1;data_in = testData6[3220];
@(posedge clk);
#1;data_in = testData6[3221];
@(posedge clk);
#1;data_in = testData6[3222];
@(posedge clk);
#1;data_in = testData6[3223];
@(posedge clk);
#1;data_in = testData6[3224];
@(posedge clk);
#1;data_in = testData6[3225];
@(posedge clk);
#1;data_in = testData6[3226];
@(posedge clk);
#1;data_in = testData6[3227];
@(posedge clk);
#1;data_in = testData6[3228];
@(posedge clk);
#1;data_in = testData6[3229];
@(posedge clk);
#1;data_in = testData6[3230];
@(posedge clk);
#1;data_in = testData6[3231];
@(posedge clk);
#1;data_in = testData6[3232];
@(posedge clk);
#1;data_in = testData6[3233];
@(posedge clk);
#1;data_in = testData6[3234];
@(posedge clk);
#1;data_in = testData6[3235];
@(posedge clk);
#1;data_in = testData6[3236];
@(posedge clk);
#1;data_in = testData6[3237];
@(posedge clk);
#1;data_in = testData6[3238];
@(posedge clk);
#1;data_in = testData6[3239];
@(posedge clk);
#1;data_in = testData6[3240];
@(posedge clk);
#1;data_in = testData6[3241];
@(posedge clk);
#1;data_in = testData6[3242];
@(posedge clk);
#1;data_in = testData6[3243];
@(posedge clk);
#1;data_in = testData6[3244];
@(posedge clk);
#1;data_in = testData6[3245];
@(posedge clk);
#1;data_in = testData6[3246];
@(posedge clk);
#1;data_in = testData6[3247];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3248]; 
@(posedge clk);
#1;data_in = testData6[3249];
@(posedge clk);
#1;data_in = testData6[3250];
@(posedge clk);
#1;data_in = testData6[3251];
@(posedge clk);
#1;data_in = testData6[3252];
@(posedge clk);
#1;data_in = testData6[3253];
@(posedge clk);
#1;data_in = testData6[3254];
@(posedge clk);
#1;data_in = testData6[3255];
@(posedge clk);
#1;data_in = testData6[3256];
@(posedge clk);
#1;data_in = testData6[3257];
@(posedge clk);
#1;data_in = testData6[3258];
@(posedge clk);
#1;data_in = testData6[3259];
@(posedge clk);
#1;data_in = testData6[3260];
@(posedge clk);
#1;data_in = testData6[3261];
@(posedge clk);
#1;data_in = testData6[3262];
@(posedge clk);
#1;data_in = testData6[3263];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3264];
@(posedge clk);
#1;data_in = testData6[3265];
@(posedge clk);
#1;data_in = testData6[3266];
@(posedge clk);
#1;data_in = testData6[3267];
@(posedge clk);
#1;data_in = testData6[3268];
@(posedge clk);
#1;data_in = testData6[3269];
@(posedge clk);
#1;data_in = testData6[3270];
@(posedge clk);
#1;data_in = testData6[3271];
@(posedge clk);
#1;data_in = testData6[3272];
@(posedge clk);
#1;data_in = testData6[3273];
@(posedge clk);
#1;data_in = testData6[3274];
@(posedge clk);
#1;data_in = testData6[3275];
@(posedge clk);
#1;data_in = testData6[3276];
@(posedge clk);
#1;data_in = testData6[3277];
@(posedge clk);
#1;data_in = testData6[3278];
@(posedge clk);
#1;data_in = testData6[3279];
@(posedge clk);
#1;data_in = testData6[3280];
@(posedge clk);
#1;data_in = testData6[3281];
@(posedge clk);
#1;data_in = testData6[3282];
@(posedge clk);
#1;data_in = testData6[3283];
@(posedge clk);
#1;data_in = testData6[3284];
@(posedge clk);
#1;data_in = testData6[3285];
@(posedge clk);
#1;data_in = testData6[3286];
@(posedge clk);
#1;data_in = testData6[3287];
@(posedge clk);
#1;data_in = testData6[3288];
@(posedge clk);
#1;data_in = testData6[3289];
@(posedge clk);
#1;data_in = testData6[3290];
@(posedge clk);
#1;data_in = testData6[3291];
@(posedge clk);
#1;data_in = testData6[3292];
@(posedge clk);
#1;data_in = testData6[3293];
@(posedge clk);
#1;data_in = testData6[3294];
@(posedge clk);
#1;data_in = testData6[3295];
@(posedge clk);
#1;data_in = testData6[3296];
@(posedge clk);
#1;data_in = testData6[3297];
@(posedge clk);
#1;data_in = testData6[3298];
@(posedge clk);
#1;data_in = testData6[3299];
@(posedge clk);
#1;data_in = testData6[3300];
@(posedge clk);
#1;data_in = testData6[3301];
@(posedge clk);
#1;data_in = testData6[3302];
@(posedge clk);
#1;data_in = testData6[3303];
@(posedge clk);
#1;data_in = testData6[3304];
@(posedge clk);
#1;data_in = testData6[3305];
@(posedge clk);
#1;data_in = testData6[3306];
@(posedge clk);
#1;data_in = testData6[3307];
@(posedge clk);
#1;data_in = testData6[3308];
@(posedge clk);
#1;data_in = testData6[3309];
@(posedge clk);
#1;data_in = testData6[3310];
@(posedge clk);
#1;data_in = testData6[3311];
@(posedge clk);
#1;data_in = testData6[3312];
@(posedge clk);
#1;data_in = testData6[3313];
@(posedge clk);
#1;data_in = testData6[3314];
@(posedge clk);
#1;data_in = testData6[3315];
@(posedge clk);
#1;data_in = testData6[3316];
@(posedge clk);
#1;data_in = testData6[3317];
@(posedge clk);
#1;data_in = testData6[3318];
@(posedge clk);
#1;data_in = testData6[3319];
@(posedge clk);
#1;data_in = testData6[3320];
@(posedge clk);
#1;data_in = testData6[3321];
@(posedge clk);
#1;data_in = testData6[3322];
@(posedge clk);
#1;data_in = testData6[3323];
@(posedge clk);
#1;data_in = testData6[3324];
@(posedge clk);
#1;data_in = testData6[3325];
@(posedge clk);
#1;data_in = testData6[3326];
@(posedge clk);
#1;data_in = testData6[3327];
@(posedge clk);
#1;data_in = testData6[3328];
@(posedge clk);
#1;data_in = testData6[3329];
@(posedge clk);
#1;data_in = testData6[3330];
@(posedge clk);
#1;data_in = testData6[3331];
@(posedge clk);
#1;data_in = testData6[3332];
@(posedge clk);
#1;data_in = testData6[3333];
@(posedge clk);
#1;data_in = testData6[3334];
@(posedge clk);
#1;data_in = testData6[3335];
@(posedge clk);
#1;data_in = testData6[3336];
@(posedge clk);
#1;data_in = testData6[3337];
@(posedge clk);
#1;data_in = testData6[3338];
@(posedge clk);
#1;data_in = testData6[3339];
@(posedge clk);
#1;data_in = testData6[3340];
@(posedge clk);
#1;data_in = testData6[3341];
@(posedge clk);
#1;data_in = testData6[3342];
@(posedge clk);
#1;data_in = testData6[3343];
@(posedge clk);
#1;data_in = testData6[3344];
@(posedge clk);
#1;data_in = testData6[3345];
@(posedge clk);
#1;data_in = testData6[3346];
@(posedge clk);
#1;data_in = testData6[3347];
@(posedge clk);
#1;data_in = testData6[3348];
@(posedge clk);
#1;data_in = testData6[3349];
@(posedge clk);
#1;data_in = testData6[3350];
@(posedge clk);
#1;data_in = testData6[3351];
@(posedge clk);
#1;data_in = testData6[3352];
@(posedge clk);
#1;data_in = testData6[3353];
@(posedge clk);
#1;data_in = testData6[3354];
@(posedge clk);
#1;data_in = testData6[3355];
@(posedge clk);
#1;data_in = testData6[3356];
@(posedge clk);
#1;data_in = testData6[3357];
@(posedge clk);
#1;data_in = testData6[3358];
@(posedge clk);
#1;data_in = testData6[3359];
@(posedge clk);
#1;data_in = testData6[3360];
@(posedge clk);
#1;data_in = testData6[3361];
@(posedge clk);
#1;data_in = testData6[3362];
@(posedge clk);
#1;data_in = testData6[3363];
@(posedge clk);
#1;data_in = testData6[3364];
@(posedge clk);
#1;data_in = testData6[3365];
@(posedge clk);
#1;data_in = testData6[3366];
@(posedge clk);
#1;data_in = testData6[3367];
@(posedge clk);
#1;data_in = testData6[3368];
@(posedge clk);
#1;data_in = testData6[3369];
@(posedge clk);
#1;data_in = testData6[3370];
@(posedge clk);
#1;data_in = testData6[3371];
@(posedge clk);
#1;data_in = testData6[3372];
@(posedge clk);
#1;data_in = testData6[3373];
@(posedge clk);
#1;data_in = testData6[3374];
@(posedge clk);
#1;data_in = testData6[3375];
@(posedge clk);
#1;data_in = testData6[3376];
@(posedge clk);
#1;data_in = testData6[3377];
@(posedge clk);
#1;data_in = testData6[3378];
@(posedge clk);
#1;data_in = testData6[3379];
@(posedge clk);
#1;data_in = testData6[3380];
@(posedge clk);
#1;data_in = testData6[3381];
@(posedge clk);
#1;data_in = testData6[3382];
@(posedge clk);
#1;data_in = testData6[3383];
@(posedge clk);
#1;data_in = testData6[3384];
@(posedge clk);
#1;data_in = testData6[3385];
@(posedge clk);
#1;data_in = testData6[3386];
@(posedge clk);
#1;data_in = testData6[3387];
@(posedge clk);
#1;data_in = testData6[3388];
@(posedge clk);
#1;data_in = testData6[3389];
@(posedge clk);
#1;data_in = testData6[3390];
@(posedge clk);
#1;data_in = testData6[3391];
@(posedge clk);
#1;data_in = testData6[3392];
@(posedge clk);
#1;data_in = testData6[3393];
@(posedge clk);
#1;data_in = testData6[3394];
@(posedge clk);
#1;data_in = testData6[3395];
@(posedge clk);
#1;data_in = testData6[3396];
@(posedge clk);
#1;data_in = testData6[3397];
@(posedge clk);
#1;data_in = testData6[3398];
@(posedge clk);
#1;data_in = testData6[3399];
@(posedge clk);
#1;data_in = testData6[3400];
@(posedge clk);
#1;data_in = testData6[3401];
@(posedge clk);
#1;data_in = testData6[3402];
@(posedge clk);
#1;data_in = testData6[3403];
@(posedge clk);
#1;data_in = testData6[3404];
@(posedge clk);
#1;data_in = testData6[3405];
@(posedge clk);
#1;data_in = testData6[3406];
@(posedge clk);
#1;data_in = testData6[3407];
@(posedge clk);
#1;data_in = testData6[3408];
@(posedge clk);
#1;data_in = testData6[3409];
@(posedge clk);
#1;data_in = testData6[3410];
@(posedge clk);
#1;data_in = testData6[3411];
@(posedge clk);
#1;data_in = testData6[3412];
@(posedge clk);
#1;data_in = testData6[3413];
@(posedge clk);
#1;data_in = testData6[3414];
@(posedge clk);
#1;data_in = testData6[3415];
@(posedge clk);
#1;data_in = testData6[3416];
@(posedge clk);
#1;data_in = testData6[3417];
@(posedge clk);
#1;data_in = testData6[3418];
@(posedge clk);
#1;data_in = testData6[3419];
@(posedge clk);
#1;data_in = testData6[3420];
@(posedge clk);
#1;data_in = testData6[3421];
@(posedge clk);
#1;data_in = testData6[3422];
@(posedge clk);
#1;data_in = testData6[3423];
@(posedge clk);
#1;data_in = testData6[3424];
@(posedge clk);
#1;data_in = testData6[3425];
@(posedge clk);
#1;data_in = testData6[3426];
@(posedge clk);
#1;data_in = testData6[3427];
@(posedge clk);
#1;data_in = testData6[3428];
@(posedge clk);
#1;data_in = testData6[3429];
@(posedge clk);
#1;data_in = testData6[3430];
@(posedge clk);
#1;data_in = testData6[3431];
@(posedge clk);
#1;data_in = testData6[3432];
@(posedge clk);
#1;data_in = testData6[3433];
@(posedge clk);
#1;data_in = testData6[3434];
@(posedge clk);
#1;data_in = testData6[3435];
@(posedge clk);
#1;data_in = testData6[3436];
@(posedge clk);
#1;data_in = testData6[3437];
@(posedge clk);
#1;data_in = testData6[3438];
@(posedge clk);
#1;data_in = testData6[3439];
@(posedge clk);
#1;data_in = testData6[3440];
@(posedge clk);
#1;data_in = testData6[3441];
@(posedge clk);
#1;data_in = testData6[3442];
@(posedge clk);
#1;data_in = testData6[3443];
@(posedge clk);
#1;data_in = testData6[3444];
@(posedge clk);
#1;data_in = testData6[3445];
@(posedge clk);
#1;data_in = testData6[3446];
@(posedge clk);
#1;data_in = testData6[3447];
@(posedge clk);
#1;data_in = testData6[3448];
@(posedge clk);
#1;data_in = testData6[3449];
@(posedge clk);
#1;data_in = testData6[3450];
@(posedge clk);
#1;data_in = testData6[3451];
@(posedge clk);
#1;data_in = testData6[3452];
@(posedge clk);
#1;data_in = testData6[3453];
@(posedge clk);
#1;data_in = testData6[3454];
@(posedge clk);
#1;data_in = testData6[3455];
@(posedge clk);
#1;data_in = testData6[3456];
@(posedge clk);
#1;data_in = testData6[3457];
@(posedge clk);
#1;data_in = testData6[3458];
@(posedge clk);
#1;data_in = testData6[3459];
@(posedge clk);
#1;data_in = testData6[3460];
@(posedge clk);
#1;data_in = testData6[3461];
@(posedge clk);
#1;data_in = testData6[3462];
@(posedge clk);
#1;data_in = testData6[3463];
@(posedge clk);
#1;data_in = testData6[3464];
@(posedge clk);
#1;data_in = testData6[3465];
@(posedge clk);
#1;data_in = testData6[3466];
@(posedge clk);
#1;data_in = testData6[3467];
@(posedge clk);
#1;data_in = testData6[3468];
@(posedge clk);
#1;data_in = testData6[3469];
@(posedge clk);
#1;data_in = testData6[3470];
@(posedge clk);
#1;data_in = testData6[3471];
@(posedge clk);
#1;data_in = testData6[3472];
@(posedge clk);
#1;data_in = testData6[3473];
@(posedge clk);
#1;data_in = testData6[3474];
@(posedge clk);
#1;data_in = testData6[3475];
@(posedge clk);
#1;data_in = testData6[3476];
@(posedge clk);
#1;data_in = testData6[3477];
@(posedge clk);
#1;data_in = testData6[3478];
@(posedge clk);
#1;data_in = testData6[3479];
@(posedge clk);
#1;data_in = testData6[3480];
@(posedge clk);
#1;data_in = testData6[3481];
@(posedge clk);
#1;data_in = testData6[3482];
@(posedge clk);
#1;data_in = testData6[3483];
@(posedge clk);
#1;data_in = testData6[3484];
@(posedge clk);
#1;data_in = testData6[3485];
@(posedge clk);
#1;data_in = testData6[3486];
@(posedge clk);
#1;data_in = testData6[3487];
@(posedge clk);
#1;data_in = testData6[3488];
@(posedge clk);
#1;data_in = testData6[3489];
@(posedge clk);
#1;data_in = testData6[3490];
@(posedge clk);
#1;data_in = testData6[3491];
@(posedge clk);
#1;data_in = testData6[3492];
@(posedge clk);
#1;data_in = testData6[3493];
@(posedge clk);
#1;data_in = testData6[3494];
@(posedge clk);
#1;data_in = testData6[3495];
@(posedge clk);
#1;data_in = testData6[3496];
@(posedge clk);
#1;data_in = testData6[3497];
@(posedge clk);
#1;data_in = testData6[3498];
@(posedge clk);
#1;data_in = testData6[3499];
@(posedge clk);
#1;data_in = testData6[3500];
@(posedge clk);
#1;data_in = testData6[3501];
@(posedge clk);
#1;data_in = testData6[3502];
@(posedge clk);
#1;data_in = testData6[3503];
@(posedge clk);
#1;data_in = testData6[3504];
@(posedge clk);
#1;data_in = testData6[3505];
@(posedge clk);
#1;data_in = testData6[3506];
@(posedge clk);
#1;data_in = testData6[3507];
@(posedge clk);
#1;data_in = testData6[3508];
@(posedge clk);
#1;data_in = testData6[3509];
@(posedge clk);
#1;data_in = testData6[3510];
@(posedge clk);
#1;data_in = testData6[3511];
@(posedge clk);
#1;data_in = testData6[3512];
@(posedge clk);
#1;data_in = testData6[3513];
@(posedge clk);
#1;data_in = testData6[3514];
@(posedge clk);
#1;data_in = testData6[3515];
@(posedge clk);
#1;data_in = testData6[3516];
@(posedge clk);
#1;data_in = testData6[3517];
@(posedge clk);
#1;data_in = testData6[3518];
@(posedge clk);
#1;data_in = testData6[3519];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3520]; 
@(posedge clk);
#1;data_in = testData6[3521];
@(posedge clk);
#1;data_in = testData6[3522];
@(posedge clk);
#1;data_in = testData6[3523];
@(posedge clk);
#1;data_in = testData6[3524];
@(posedge clk);
#1;data_in = testData6[3525];
@(posedge clk);
#1;data_in = testData6[3526];
@(posedge clk);
#1;data_in = testData6[3527];
@(posedge clk);
#1;data_in = testData6[3528];
@(posedge clk);
#1;data_in = testData6[3529];
@(posedge clk);
#1;data_in = testData6[3530];
@(posedge clk);
#1;data_in = testData6[3531];
@(posedge clk);
#1;data_in = testData6[3532];
@(posedge clk);
#1;data_in = testData6[3533];
@(posedge clk);
#1;data_in = testData6[3534];
@(posedge clk);
#1;data_in = testData6[3535];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3536];
@(posedge clk);
#1;data_in = testData6[3537];
@(posedge clk);
#1;data_in = testData6[3538];
@(posedge clk);
#1;data_in = testData6[3539];
@(posedge clk);
#1;data_in = testData6[3540];
@(posedge clk);
#1;data_in = testData6[3541];
@(posedge clk);
#1;data_in = testData6[3542];
@(posedge clk);
#1;data_in = testData6[3543];
@(posedge clk);
#1;data_in = testData6[3544];
@(posedge clk);
#1;data_in = testData6[3545];
@(posedge clk);
#1;data_in = testData6[3546];
@(posedge clk);
#1;data_in = testData6[3547];
@(posedge clk);
#1;data_in = testData6[3548];
@(posedge clk);
#1;data_in = testData6[3549];
@(posedge clk);
#1;data_in = testData6[3550];
@(posedge clk);
#1;data_in = testData6[3551];
@(posedge clk);
#1;data_in = testData6[3552];
@(posedge clk);
#1;data_in = testData6[3553];
@(posedge clk);
#1;data_in = testData6[3554];
@(posedge clk);
#1;data_in = testData6[3555];
@(posedge clk);
#1;data_in = testData6[3556];
@(posedge clk);
#1;data_in = testData6[3557];
@(posedge clk);
#1;data_in = testData6[3558];
@(posedge clk);
#1;data_in = testData6[3559];
@(posedge clk);
#1;data_in = testData6[3560];
@(posedge clk);
#1;data_in = testData6[3561];
@(posedge clk);
#1;data_in = testData6[3562];
@(posedge clk);
#1;data_in = testData6[3563];
@(posedge clk);
#1;data_in = testData6[3564];
@(posedge clk);
#1;data_in = testData6[3565];
@(posedge clk);
#1;data_in = testData6[3566];
@(posedge clk);
#1;data_in = testData6[3567];
@(posedge clk);
#1;data_in = testData6[3568];
@(posedge clk);
#1;data_in = testData6[3569];
@(posedge clk);
#1;data_in = testData6[3570];
@(posedge clk);
#1;data_in = testData6[3571];
@(posedge clk);
#1;data_in = testData6[3572];
@(posedge clk);
#1;data_in = testData6[3573];
@(posedge clk);
#1;data_in = testData6[3574];
@(posedge clk);
#1;data_in = testData6[3575];
@(posedge clk);
#1;data_in = testData6[3576];
@(posedge clk);
#1;data_in = testData6[3577];
@(posedge clk);
#1;data_in = testData6[3578];
@(posedge clk);
#1;data_in = testData6[3579];
@(posedge clk);
#1;data_in = testData6[3580];
@(posedge clk);
#1;data_in = testData6[3581];
@(posedge clk);
#1;data_in = testData6[3582];
@(posedge clk);
#1;data_in = testData6[3583];
@(posedge clk);
#1;data_in = testData6[3584];
@(posedge clk);
#1;data_in = testData6[3585];
@(posedge clk);
#1;data_in = testData6[3586];
@(posedge clk);
#1;data_in = testData6[3587];
@(posedge clk);
#1;data_in = testData6[3588];
@(posedge clk);
#1;data_in = testData6[3589];
@(posedge clk);
#1;data_in = testData6[3590];
@(posedge clk);
#1;data_in = testData6[3591];
@(posedge clk);
#1;data_in = testData6[3592];
@(posedge clk);
#1;data_in = testData6[3593];
@(posedge clk);
#1;data_in = testData6[3594];
@(posedge clk);
#1;data_in = testData6[3595];
@(posedge clk);
#1;data_in = testData6[3596];
@(posedge clk);
#1;data_in = testData6[3597];
@(posedge clk);
#1;data_in = testData6[3598];
@(posedge clk);
#1;data_in = testData6[3599];
@(posedge clk);
#1;data_in = testData6[3600];
@(posedge clk);
#1;data_in = testData6[3601];
@(posedge clk);
#1;data_in = testData6[3602];
@(posedge clk);
#1;data_in = testData6[3603];
@(posedge clk);
#1;data_in = testData6[3604];
@(posedge clk);
#1;data_in = testData6[3605];
@(posedge clk);
#1;data_in = testData6[3606];
@(posedge clk);
#1;data_in = testData6[3607];
@(posedge clk);
#1;data_in = testData6[3608];
@(posedge clk);
#1;data_in = testData6[3609];
@(posedge clk);
#1;data_in = testData6[3610];
@(posedge clk);
#1;data_in = testData6[3611];
@(posedge clk);
#1;data_in = testData6[3612];
@(posedge clk);
#1;data_in = testData6[3613];
@(posedge clk);
#1;data_in = testData6[3614];
@(posedge clk);
#1;data_in = testData6[3615];
@(posedge clk);
#1;data_in = testData6[3616];
@(posedge clk);
#1;data_in = testData6[3617];
@(posedge clk);
#1;data_in = testData6[3618];
@(posedge clk);
#1;data_in = testData6[3619];
@(posedge clk);
#1;data_in = testData6[3620];
@(posedge clk);
#1;data_in = testData6[3621];
@(posedge clk);
#1;data_in = testData6[3622];
@(posedge clk);
#1;data_in = testData6[3623];
@(posedge clk);
#1;data_in = testData6[3624];
@(posedge clk);
#1;data_in = testData6[3625];
@(posedge clk);
#1;data_in = testData6[3626];
@(posedge clk);
#1;data_in = testData6[3627];
@(posedge clk);
#1;data_in = testData6[3628];
@(posedge clk);
#1;data_in = testData6[3629];
@(posedge clk);
#1;data_in = testData6[3630];
@(posedge clk);
#1;data_in = testData6[3631];
@(posedge clk);
#1;data_in = testData6[3632];
@(posedge clk);
#1;data_in = testData6[3633];
@(posedge clk);
#1;data_in = testData6[3634];
@(posedge clk);
#1;data_in = testData6[3635];
@(posedge clk);
#1;data_in = testData6[3636];
@(posedge clk);
#1;data_in = testData6[3637];
@(posedge clk);
#1;data_in = testData6[3638];
@(posedge clk);
#1;data_in = testData6[3639];
@(posedge clk);
#1;data_in = testData6[3640];
@(posedge clk);
#1;data_in = testData6[3641];
@(posedge clk);
#1;data_in = testData6[3642];
@(posedge clk);
#1;data_in = testData6[3643];
@(posedge clk);
#1;data_in = testData6[3644];
@(posedge clk);
#1;data_in = testData6[3645];
@(posedge clk);
#1;data_in = testData6[3646];
@(posedge clk);
#1;data_in = testData6[3647];
@(posedge clk);
#1;data_in = testData6[3648];
@(posedge clk);
#1;data_in = testData6[3649];
@(posedge clk);
#1;data_in = testData6[3650];
@(posedge clk);
#1;data_in = testData6[3651];
@(posedge clk);
#1;data_in = testData6[3652];
@(posedge clk);
#1;data_in = testData6[3653];
@(posedge clk);
#1;data_in = testData6[3654];
@(posedge clk);
#1;data_in = testData6[3655];
@(posedge clk);
#1;data_in = testData6[3656];
@(posedge clk);
#1;data_in = testData6[3657];
@(posedge clk);
#1;data_in = testData6[3658];
@(posedge clk);
#1;data_in = testData6[3659];
@(posedge clk);
#1;data_in = testData6[3660];
@(posedge clk);
#1;data_in = testData6[3661];
@(posedge clk);
#1;data_in = testData6[3662];
@(posedge clk);
#1;data_in = testData6[3663];
@(posedge clk);
#1;data_in = testData6[3664];
@(posedge clk);
#1;data_in = testData6[3665];
@(posedge clk);
#1;data_in = testData6[3666];
@(posedge clk);
#1;data_in = testData6[3667];
@(posedge clk);
#1;data_in = testData6[3668];
@(posedge clk);
#1;data_in = testData6[3669];
@(posedge clk);
#1;data_in = testData6[3670];
@(posedge clk);
#1;data_in = testData6[3671];
@(posedge clk);
#1;data_in = testData6[3672];
@(posedge clk);
#1;data_in = testData6[3673];
@(posedge clk);
#1;data_in = testData6[3674];
@(posedge clk);
#1;data_in = testData6[3675];
@(posedge clk);
#1;data_in = testData6[3676];
@(posedge clk);
#1;data_in = testData6[3677];
@(posedge clk);
#1;data_in = testData6[3678];
@(posedge clk);
#1;data_in = testData6[3679];
@(posedge clk);
#1;data_in = testData6[3680];
@(posedge clk);
#1;data_in = testData6[3681];
@(posedge clk);
#1;data_in = testData6[3682];
@(posedge clk);
#1;data_in = testData6[3683];
@(posedge clk);
#1;data_in = testData6[3684];
@(posedge clk);
#1;data_in = testData6[3685];
@(posedge clk);
#1;data_in = testData6[3686];
@(posedge clk);
#1;data_in = testData6[3687];
@(posedge clk);
#1;data_in = testData6[3688];
@(posedge clk);
#1;data_in = testData6[3689];
@(posedge clk);
#1;data_in = testData6[3690];
@(posedge clk);
#1;data_in = testData6[3691];
@(posedge clk);
#1;data_in = testData6[3692];
@(posedge clk);
#1;data_in = testData6[3693];
@(posedge clk);
#1;data_in = testData6[3694];
@(posedge clk);
#1;data_in = testData6[3695];
@(posedge clk);
#1;data_in = testData6[3696];
@(posedge clk);
#1;data_in = testData6[3697];
@(posedge clk);
#1;data_in = testData6[3698];
@(posedge clk);
#1;data_in = testData6[3699];
@(posedge clk);
#1;data_in = testData6[3700];
@(posedge clk);
#1;data_in = testData6[3701];
@(posedge clk);
#1;data_in = testData6[3702];
@(posedge clk);
#1;data_in = testData6[3703];
@(posedge clk);
#1;data_in = testData6[3704];
@(posedge clk);
#1;data_in = testData6[3705];
@(posedge clk);
#1;data_in = testData6[3706];
@(posedge clk);
#1;data_in = testData6[3707];
@(posedge clk);
#1;data_in = testData6[3708];
@(posedge clk);
#1;data_in = testData6[3709];
@(posedge clk);
#1;data_in = testData6[3710];
@(posedge clk);
#1;data_in = testData6[3711];
@(posedge clk);
#1;data_in = testData6[3712];
@(posedge clk);
#1;data_in = testData6[3713];
@(posedge clk);
#1;data_in = testData6[3714];
@(posedge clk);
#1;data_in = testData6[3715];
@(posedge clk);
#1;data_in = testData6[3716];
@(posedge clk);
#1;data_in = testData6[3717];
@(posedge clk);
#1;data_in = testData6[3718];
@(posedge clk);
#1;data_in = testData6[3719];
@(posedge clk);
#1;data_in = testData6[3720];
@(posedge clk);
#1;data_in = testData6[3721];
@(posedge clk);
#1;data_in = testData6[3722];
@(posedge clk);
#1;data_in = testData6[3723];
@(posedge clk);
#1;data_in = testData6[3724];
@(posedge clk);
#1;data_in = testData6[3725];
@(posedge clk);
#1;data_in = testData6[3726];
@(posedge clk);
#1;data_in = testData6[3727];
@(posedge clk);
#1;data_in = testData6[3728];
@(posedge clk);
#1;data_in = testData6[3729];
@(posedge clk);
#1;data_in = testData6[3730];
@(posedge clk);
#1;data_in = testData6[3731];
@(posedge clk);
#1;data_in = testData6[3732];
@(posedge clk);
#1;data_in = testData6[3733];
@(posedge clk);
#1;data_in = testData6[3734];
@(posedge clk);
#1;data_in = testData6[3735];
@(posedge clk);
#1;data_in = testData6[3736];
@(posedge clk);
#1;data_in = testData6[3737];
@(posedge clk);
#1;data_in = testData6[3738];
@(posedge clk);
#1;data_in = testData6[3739];
@(posedge clk);
#1;data_in = testData6[3740];
@(posedge clk);
#1;data_in = testData6[3741];
@(posedge clk);
#1;data_in = testData6[3742];
@(posedge clk);
#1;data_in = testData6[3743];
@(posedge clk);
#1;data_in = testData6[3744];
@(posedge clk);
#1;data_in = testData6[3745];
@(posedge clk);
#1;data_in = testData6[3746];
@(posedge clk);
#1;data_in = testData6[3747];
@(posedge clk);
#1;data_in = testData6[3748];
@(posedge clk);
#1;data_in = testData6[3749];
@(posedge clk);
#1;data_in = testData6[3750];
@(posedge clk);
#1;data_in = testData6[3751];
@(posedge clk);
#1;data_in = testData6[3752];
@(posedge clk);
#1;data_in = testData6[3753];
@(posedge clk);
#1;data_in = testData6[3754];
@(posedge clk);
#1;data_in = testData6[3755];
@(posedge clk);
#1;data_in = testData6[3756];
@(posedge clk);
#1;data_in = testData6[3757];
@(posedge clk);
#1;data_in = testData6[3758];
@(posedge clk);
#1;data_in = testData6[3759];
@(posedge clk);
#1;data_in = testData6[3760];
@(posedge clk);
#1;data_in = testData6[3761];
@(posedge clk);
#1;data_in = testData6[3762];
@(posedge clk);
#1;data_in = testData6[3763];
@(posedge clk);
#1;data_in = testData6[3764];
@(posedge clk);
#1;data_in = testData6[3765];
@(posedge clk);
#1;data_in = testData6[3766];
@(posedge clk);
#1;data_in = testData6[3767];
@(posedge clk);
#1;data_in = testData6[3768];
@(posedge clk);
#1;data_in = testData6[3769];
@(posedge clk);
#1;data_in = testData6[3770];
@(posedge clk);
#1;data_in = testData6[3771];
@(posedge clk);
#1;data_in = testData6[3772];
@(posedge clk);
#1;data_in = testData6[3773];
@(posedge clk);
#1;data_in = testData6[3774];
@(posedge clk);
#1;data_in = testData6[3775];
@(posedge clk);
#1;data_in = testData6[3776];
@(posedge clk);
#1;data_in = testData6[3777];
@(posedge clk);
#1;data_in = testData6[3778];
@(posedge clk);
#1;data_in = testData6[3779];
@(posedge clk);
#1;data_in = testData6[3780];
@(posedge clk);
#1;data_in = testData6[3781];
@(posedge clk);
#1;data_in = testData6[3782];
@(posedge clk);
#1;data_in = testData6[3783];
@(posedge clk);
#1;data_in = testData6[3784];
@(posedge clk);
#1;data_in = testData6[3785];
@(posedge clk);
#1;data_in = testData6[3786];
@(posedge clk);
#1;data_in = testData6[3787];
@(posedge clk);
#1;data_in = testData6[3788];
@(posedge clk);
#1;data_in = testData6[3789];
@(posedge clk);
#1;data_in = testData6[3790];
@(posedge clk);
#1;data_in = testData6[3791];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3792]; 
@(posedge clk);
#1;data_in = testData6[3793];
@(posedge clk);
#1;data_in = testData6[3794];
@(posedge clk);
#1;data_in = testData6[3795];
@(posedge clk);
#1;data_in = testData6[3796];
@(posedge clk);
#1;data_in = testData6[3797];
@(posedge clk);
#1;data_in = testData6[3798];
@(posedge clk);
#1;data_in = testData6[3799];
@(posedge clk);
#1;data_in = testData6[3800];
@(posedge clk);
#1;data_in = testData6[3801];
@(posedge clk);
#1;data_in = testData6[3802];
@(posedge clk);
#1;data_in = testData6[3803];
@(posedge clk);
#1;data_in = testData6[3804];
@(posedge clk);
#1;data_in = testData6[3805];
@(posedge clk);
#1;data_in = testData6[3806];
@(posedge clk);
#1;data_in = testData6[3807];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3808];
@(posedge clk);
#1;data_in = testData6[3809];
@(posedge clk);
#1;data_in = testData6[3810];
@(posedge clk);
#1;data_in = testData6[3811];
@(posedge clk);
#1;data_in = testData6[3812];
@(posedge clk);
#1;data_in = testData6[3813];
@(posedge clk);
#1;data_in = testData6[3814];
@(posedge clk);
#1;data_in = testData6[3815];
@(posedge clk);
#1;data_in = testData6[3816];
@(posedge clk);
#1;data_in = testData6[3817];
@(posedge clk);
#1;data_in = testData6[3818];
@(posedge clk);
#1;data_in = testData6[3819];
@(posedge clk);
#1;data_in = testData6[3820];
@(posedge clk);
#1;data_in = testData6[3821];
@(posedge clk);
#1;data_in = testData6[3822];
@(posedge clk);
#1;data_in = testData6[3823];
@(posedge clk);
#1;data_in = testData6[3824];
@(posedge clk);
#1;data_in = testData6[3825];
@(posedge clk);
#1;data_in = testData6[3826];
@(posedge clk);
#1;data_in = testData6[3827];
@(posedge clk);
#1;data_in = testData6[3828];
@(posedge clk);
#1;data_in = testData6[3829];
@(posedge clk);
#1;data_in = testData6[3830];
@(posedge clk);
#1;data_in = testData6[3831];
@(posedge clk);
#1;data_in = testData6[3832];
@(posedge clk);
#1;data_in = testData6[3833];
@(posedge clk);
#1;data_in = testData6[3834];
@(posedge clk);
#1;data_in = testData6[3835];
@(posedge clk);
#1;data_in = testData6[3836];
@(posedge clk);
#1;data_in = testData6[3837];
@(posedge clk);
#1;data_in = testData6[3838];
@(posedge clk);
#1;data_in = testData6[3839];
@(posedge clk);
#1;data_in = testData6[3840];
@(posedge clk);
#1;data_in = testData6[3841];
@(posedge clk);
#1;data_in = testData6[3842];
@(posedge clk);
#1;data_in = testData6[3843];
@(posedge clk);
#1;data_in = testData6[3844];
@(posedge clk);
#1;data_in = testData6[3845];
@(posedge clk);
#1;data_in = testData6[3846];
@(posedge clk);
#1;data_in = testData6[3847];
@(posedge clk);
#1;data_in = testData6[3848];
@(posedge clk);
#1;data_in = testData6[3849];
@(posedge clk);
#1;data_in = testData6[3850];
@(posedge clk);
#1;data_in = testData6[3851];
@(posedge clk);
#1;data_in = testData6[3852];
@(posedge clk);
#1;data_in = testData6[3853];
@(posedge clk);
#1;data_in = testData6[3854];
@(posedge clk);
#1;data_in = testData6[3855];
@(posedge clk);
#1;data_in = testData6[3856];
@(posedge clk);
#1;data_in = testData6[3857];
@(posedge clk);
#1;data_in = testData6[3858];
@(posedge clk);
#1;data_in = testData6[3859];
@(posedge clk);
#1;data_in = testData6[3860];
@(posedge clk);
#1;data_in = testData6[3861];
@(posedge clk);
#1;data_in = testData6[3862];
@(posedge clk);
#1;data_in = testData6[3863];
@(posedge clk);
#1;data_in = testData6[3864];
@(posedge clk);
#1;data_in = testData6[3865];
@(posedge clk);
#1;data_in = testData6[3866];
@(posedge clk);
#1;data_in = testData6[3867];
@(posedge clk);
#1;data_in = testData6[3868];
@(posedge clk);
#1;data_in = testData6[3869];
@(posedge clk);
#1;data_in = testData6[3870];
@(posedge clk);
#1;data_in = testData6[3871];
@(posedge clk);
#1;data_in = testData6[3872];
@(posedge clk);
#1;data_in = testData6[3873];
@(posedge clk);
#1;data_in = testData6[3874];
@(posedge clk);
#1;data_in = testData6[3875];
@(posedge clk);
#1;data_in = testData6[3876];
@(posedge clk);
#1;data_in = testData6[3877];
@(posedge clk);
#1;data_in = testData6[3878];
@(posedge clk);
#1;data_in = testData6[3879];
@(posedge clk);
#1;data_in = testData6[3880];
@(posedge clk);
#1;data_in = testData6[3881];
@(posedge clk);
#1;data_in = testData6[3882];
@(posedge clk);
#1;data_in = testData6[3883];
@(posedge clk);
#1;data_in = testData6[3884];
@(posedge clk);
#1;data_in = testData6[3885];
@(posedge clk);
#1;data_in = testData6[3886];
@(posedge clk);
#1;data_in = testData6[3887];
@(posedge clk);
#1;data_in = testData6[3888];
@(posedge clk);
#1;data_in = testData6[3889];
@(posedge clk);
#1;data_in = testData6[3890];
@(posedge clk);
#1;data_in = testData6[3891];
@(posedge clk);
#1;data_in = testData6[3892];
@(posedge clk);
#1;data_in = testData6[3893];
@(posedge clk);
#1;data_in = testData6[3894];
@(posedge clk);
#1;data_in = testData6[3895];
@(posedge clk);
#1;data_in = testData6[3896];
@(posedge clk);
#1;data_in = testData6[3897];
@(posedge clk);
#1;data_in = testData6[3898];
@(posedge clk);
#1;data_in = testData6[3899];
@(posedge clk);
#1;data_in = testData6[3900];
@(posedge clk);
#1;data_in = testData6[3901];
@(posedge clk);
#1;data_in = testData6[3902];
@(posedge clk);
#1;data_in = testData6[3903];
@(posedge clk);
#1;data_in = testData6[3904];
@(posedge clk);
#1;data_in = testData6[3905];
@(posedge clk);
#1;data_in = testData6[3906];
@(posedge clk);
#1;data_in = testData6[3907];
@(posedge clk);
#1;data_in = testData6[3908];
@(posedge clk);
#1;data_in = testData6[3909];
@(posedge clk);
#1;data_in = testData6[3910];
@(posedge clk);
#1;data_in = testData6[3911];
@(posedge clk);
#1;data_in = testData6[3912];
@(posedge clk);
#1;data_in = testData6[3913];
@(posedge clk);
#1;data_in = testData6[3914];
@(posedge clk);
#1;data_in = testData6[3915];
@(posedge clk);
#1;data_in = testData6[3916];
@(posedge clk);
#1;data_in = testData6[3917];
@(posedge clk);
#1;data_in = testData6[3918];
@(posedge clk);
#1;data_in = testData6[3919];
@(posedge clk);
#1;data_in = testData6[3920];
@(posedge clk);
#1;data_in = testData6[3921];
@(posedge clk);
#1;data_in = testData6[3922];
@(posedge clk);
#1;data_in = testData6[3923];
@(posedge clk);
#1;data_in = testData6[3924];
@(posedge clk);
#1;data_in = testData6[3925];
@(posedge clk);
#1;data_in = testData6[3926];
@(posedge clk);
#1;data_in = testData6[3927];
@(posedge clk);
#1;data_in = testData6[3928];
@(posedge clk);
#1;data_in = testData6[3929];
@(posedge clk);
#1;data_in = testData6[3930];
@(posedge clk);
#1;data_in = testData6[3931];
@(posedge clk);
#1;data_in = testData6[3932];
@(posedge clk);
#1;data_in = testData6[3933];
@(posedge clk);
#1;data_in = testData6[3934];
@(posedge clk);
#1;data_in = testData6[3935];
@(posedge clk);
#1;data_in = testData6[3936];
@(posedge clk);
#1;data_in = testData6[3937];
@(posedge clk);
#1;data_in = testData6[3938];
@(posedge clk);
#1;data_in = testData6[3939];
@(posedge clk);
#1;data_in = testData6[3940];
@(posedge clk);
#1;data_in = testData6[3941];
@(posedge clk);
#1;data_in = testData6[3942];
@(posedge clk);
#1;data_in = testData6[3943];
@(posedge clk);
#1;data_in = testData6[3944];
@(posedge clk);
#1;data_in = testData6[3945];
@(posedge clk);
#1;data_in = testData6[3946];
@(posedge clk);
#1;data_in = testData6[3947];
@(posedge clk);
#1;data_in = testData6[3948];
@(posedge clk);
#1;data_in = testData6[3949];
@(posedge clk);
#1;data_in = testData6[3950];
@(posedge clk);
#1;data_in = testData6[3951];
@(posedge clk);
#1;data_in = testData6[3952];
@(posedge clk);
#1;data_in = testData6[3953];
@(posedge clk);
#1;data_in = testData6[3954];
@(posedge clk);
#1;data_in = testData6[3955];
@(posedge clk);
#1;data_in = testData6[3956];
@(posedge clk);
#1;data_in = testData6[3957];
@(posedge clk);
#1;data_in = testData6[3958];
@(posedge clk);
#1;data_in = testData6[3959];
@(posedge clk);
#1;data_in = testData6[3960];
@(posedge clk);
#1;data_in = testData6[3961];
@(posedge clk);
#1;data_in = testData6[3962];
@(posedge clk);
#1;data_in = testData6[3963];
@(posedge clk);
#1;data_in = testData6[3964];
@(posedge clk);
#1;data_in = testData6[3965];
@(posedge clk);
#1;data_in = testData6[3966];
@(posedge clk);
#1;data_in = testData6[3967];
@(posedge clk);
#1;data_in = testData6[3968];
@(posedge clk);
#1;data_in = testData6[3969];
@(posedge clk);
#1;data_in = testData6[3970];
@(posedge clk);
#1;data_in = testData6[3971];
@(posedge clk);
#1;data_in = testData6[3972];
@(posedge clk);
#1;data_in = testData6[3973];
@(posedge clk);
#1;data_in = testData6[3974];
@(posedge clk);
#1;data_in = testData6[3975];
@(posedge clk);
#1;data_in = testData6[3976];
@(posedge clk);
#1;data_in = testData6[3977];
@(posedge clk);
#1;data_in = testData6[3978];
@(posedge clk);
#1;data_in = testData6[3979];
@(posedge clk);
#1;data_in = testData6[3980];
@(posedge clk);
#1;data_in = testData6[3981];
@(posedge clk);
#1;data_in = testData6[3982];
@(posedge clk);
#1;data_in = testData6[3983];
@(posedge clk);
#1;data_in = testData6[3984];
@(posedge clk);
#1;data_in = testData6[3985];
@(posedge clk);
#1;data_in = testData6[3986];
@(posedge clk);
#1;data_in = testData6[3987];
@(posedge clk);
#1;data_in = testData6[3988];
@(posedge clk);
#1;data_in = testData6[3989];
@(posedge clk);
#1;data_in = testData6[3990];
@(posedge clk);
#1;data_in = testData6[3991];
@(posedge clk);
#1;data_in = testData6[3992];
@(posedge clk);
#1;data_in = testData6[3993];
@(posedge clk);
#1;data_in = testData6[3994];
@(posedge clk);
#1;data_in = testData6[3995];
@(posedge clk);
#1;data_in = testData6[3996];
@(posedge clk);
#1;data_in = testData6[3997];
@(posedge clk);
#1;data_in = testData6[3998];
@(posedge clk);
#1;data_in = testData6[3999];
@(posedge clk);
#1;data_in = testData6[4000];
@(posedge clk);
#1;data_in = testData6[4001];
@(posedge clk);
#1;data_in = testData6[4002];
@(posedge clk);
#1;data_in = testData6[4003];
@(posedge clk);
#1;data_in = testData6[4004];
@(posedge clk);
#1;data_in = testData6[4005];
@(posedge clk);
#1;data_in = testData6[4006];
@(posedge clk);
#1;data_in = testData6[4007];
@(posedge clk);
#1;data_in = testData6[4008];
@(posedge clk);
#1;data_in = testData6[4009];
@(posedge clk);
#1;data_in = testData6[4010];
@(posedge clk);
#1;data_in = testData6[4011];
@(posedge clk);
#1;data_in = testData6[4012];
@(posedge clk);
#1;data_in = testData6[4013];
@(posedge clk);
#1;data_in = testData6[4014];
@(posedge clk);
#1;data_in = testData6[4015];
@(posedge clk);
#1;data_in = testData6[4016];
@(posedge clk);
#1;data_in = testData6[4017];
@(posedge clk);
#1;data_in = testData6[4018];
@(posedge clk);
#1;data_in = testData6[4019];
@(posedge clk);
#1;data_in = testData6[4020];
@(posedge clk);
#1;data_in = testData6[4021];
@(posedge clk);
#1;data_in = testData6[4022];
@(posedge clk);
#1;data_in = testData6[4023];
@(posedge clk);
#1;data_in = testData6[4024];
@(posedge clk);
#1;data_in = testData6[4025];
@(posedge clk);
#1;data_in = testData6[4026];
@(posedge clk);
#1;data_in = testData6[4027];
@(posedge clk);
#1;data_in = testData6[4028];
@(posedge clk);
#1;data_in = testData6[4029];
@(posedge clk);
#1;data_in = testData6[4030];
@(posedge clk);
#1;data_in = testData6[4031];
@(posedge clk);
#1;data_in = testData6[4032];
@(posedge clk);
#1;data_in = testData6[4033];
@(posedge clk);
#1;data_in = testData6[4034];
@(posedge clk);
#1;data_in = testData6[4035];
@(posedge clk);
#1;data_in = testData6[4036];
@(posedge clk);
#1;data_in = testData6[4037];
@(posedge clk);
#1;data_in = testData6[4038];
@(posedge clk);
#1;data_in = testData6[4039];
@(posedge clk);
#1;data_in = testData6[4040];
@(posedge clk);
#1;data_in = testData6[4041];
@(posedge clk);
#1;data_in = testData6[4042];
@(posedge clk);
#1;data_in = testData6[4043];
@(posedge clk);
#1;data_in = testData6[4044];
@(posedge clk);
#1;data_in = testData6[4045];
@(posedge clk);
#1;data_in = testData6[4046];
@(posedge clk);
#1;data_in = testData6[4047];
@(posedge clk);
#1;data_in = testData6[4048];
@(posedge clk);
#1;data_in = testData6[4049];
@(posedge clk);
#1;data_in = testData6[4050];
@(posedge clk);
#1;data_in = testData6[4051];
@(posedge clk);
#1;data_in = testData6[4052];
@(posedge clk);
#1;data_in = testData6[4053];
@(posedge clk);
#1;data_in = testData6[4054];
@(posedge clk);
#1;data_in = testData6[4055];
@(posedge clk);
#1;data_in = testData6[4056];
@(posedge clk);
#1;data_in = testData6[4057];
@(posedge clk);
#1;data_in = testData6[4058];
@(posedge clk);
#1;data_in = testData6[4059];
@(posedge clk);
#1;data_in = testData6[4060];
@(posedge clk);
#1;data_in = testData6[4061];
@(posedge clk);
#1;data_in = testData6[4062];
@(posedge clk);
#1;data_in = testData6[4063];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[4064]; 
@(posedge clk);
#1;data_in = testData6[4065];
@(posedge clk);
#1;data_in = testData6[4066];
@(posedge clk);
#1;data_in = testData6[4067];
@(posedge clk);
#1;data_in = testData6[4068];
@(posedge clk);
#1;data_in = testData6[4069];
@(posedge clk);
#1;data_in = testData6[4070];
@(posedge clk);
#1;data_in = testData6[4071];
@(posedge clk);
#1;data_in = testData6[4072];
@(posedge clk);
#1;data_in = testData6[4073];
@(posedge clk);
#1;data_in = testData6[4074];
@(posedge clk);
#1;data_in = testData6[4075];
@(posedge clk);
#1;data_in = testData6[4076];
@(posedge clk);
#1;data_in = testData6[4077];
@(posedge clk);
#1;data_in = testData6[4078];
@(posedge clk);
#1;data_in = testData6[4079];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[4080];
@(posedge clk);
#1;data_in = testData6[4081];
@(posedge clk);
#1;data_in = testData6[4082];
@(posedge clk);
#1;data_in = testData6[4083];
@(posedge clk);
#1;data_in = testData6[4084];
@(posedge clk);
#1;data_in = testData6[4085];
@(posedge clk);
#1;data_in = testData6[4086];
@(posedge clk);
#1;data_in = testData6[4087];
@(posedge clk);
#1;data_in = testData6[4088];
@(posedge clk);
#1;data_in = testData6[4089];
@(posedge clk);
#1;data_in = testData6[4090];
@(posedge clk);
#1;data_in = testData6[4091];
@(posedge clk);
#1;data_in = testData6[4092];
@(posedge clk);
#1;data_in = testData6[4093];
@(posedge clk);
#1;data_in = testData6[4094];
@(posedge clk);
#1;data_in = testData6[4095];
@(posedge clk);
#1;data_in = testData6[4096];
@(posedge clk);
#1;data_in = testData6[4097];
@(posedge clk);
#1;data_in = testData6[4098];
@(posedge clk);
#1;data_in = testData6[4099];
@(posedge clk);
#1;data_in = testData6[4100];
@(posedge clk);
#1;data_in = testData6[4101];
@(posedge clk);
#1;data_in = testData6[4102];
@(posedge clk);
#1;data_in = testData6[4103];
@(posedge clk);
#1;data_in = testData6[4104];
@(posedge clk);
#1;data_in = testData6[4105];
@(posedge clk);
#1;data_in = testData6[4106];
@(posedge clk);
#1;data_in = testData6[4107];
@(posedge clk);
#1;data_in = testData6[4108];
@(posedge clk);
#1;data_in = testData6[4109];
@(posedge clk);
#1;data_in = testData6[4110];
@(posedge clk);
#1;data_in = testData6[4111];
@(posedge clk);
#1;data_in = testData6[4112];
@(posedge clk);
#1;data_in = testData6[4113];
@(posedge clk);
#1;data_in = testData6[4114];
@(posedge clk);
#1;data_in = testData6[4115];
@(posedge clk);
#1;data_in = testData6[4116];
@(posedge clk);
#1;data_in = testData6[4117];
@(posedge clk);
#1;data_in = testData6[4118];
@(posedge clk);
#1;data_in = testData6[4119];
@(posedge clk);
#1;data_in = testData6[4120];
@(posedge clk);
#1;data_in = testData6[4121];
@(posedge clk);
#1;data_in = testData6[4122];
@(posedge clk);
#1;data_in = testData6[4123];
@(posedge clk);
#1;data_in = testData6[4124];
@(posedge clk);
#1;data_in = testData6[4125];
@(posedge clk);
#1;data_in = testData6[4126];
@(posedge clk);
#1;data_in = testData6[4127];
@(posedge clk);
#1;data_in = testData6[4128];
@(posedge clk);
#1;data_in = testData6[4129];
@(posedge clk);
#1;data_in = testData6[4130];
@(posedge clk);
#1;data_in = testData6[4131];
@(posedge clk);
#1;data_in = testData6[4132];
@(posedge clk);
#1;data_in = testData6[4133];
@(posedge clk);
#1;data_in = testData6[4134];
@(posedge clk);
#1;data_in = testData6[4135];
@(posedge clk);
#1;data_in = testData6[4136];
@(posedge clk);
#1;data_in = testData6[4137];
@(posedge clk);
#1;data_in = testData6[4138];
@(posedge clk);
#1;data_in = testData6[4139];
@(posedge clk);
#1;data_in = testData6[4140];
@(posedge clk);
#1;data_in = testData6[4141];
@(posedge clk);
#1;data_in = testData6[4142];
@(posedge clk);
#1;data_in = testData6[4143];
@(posedge clk);
#1;data_in = testData6[4144];
@(posedge clk);
#1;data_in = testData6[4145];
@(posedge clk);
#1;data_in = testData6[4146];
@(posedge clk);
#1;data_in = testData6[4147];
@(posedge clk);
#1;data_in = testData6[4148];
@(posedge clk);
#1;data_in = testData6[4149];
@(posedge clk);
#1;data_in = testData6[4150];
@(posedge clk);
#1;data_in = testData6[4151];
@(posedge clk);
#1;data_in = testData6[4152];
@(posedge clk);
#1;data_in = testData6[4153];
@(posedge clk);
#1;data_in = testData6[4154];
@(posedge clk);
#1;data_in = testData6[4155];
@(posedge clk);
#1;data_in = testData6[4156];
@(posedge clk);
#1;data_in = testData6[4157];
@(posedge clk);
#1;data_in = testData6[4158];
@(posedge clk);
#1;data_in = testData6[4159];
@(posedge clk);
#1;data_in = testData6[4160];
@(posedge clk);
#1;data_in = testData6[4161];
@(posedge clk);
#1;data_in = testData6[4162];
@(posedge clk);
#1;data_in = testData6[4163];
@(posedge clk);
#1;data_in = testData6[4164];
@(posedge clk);
#1;data_in = testData6[4165];
@(posedge clk);
#1;data_in = testData6[4166];
@(posedge clk);
#1;data_in = testData6[4167];
@(posedge clk);
#1;data_in = testData6[4168];
@(posedge clk);
#1;data_in = testData6[4169];
@(posedge clk);
#1;data_in = testData6[4170];
@(posedge clk);
#1;data_in = testData6[4171];
@(posedge clk);
#1;data_in = testData6[4172];
@(posedge clk);
#1;data_in = testData6[4173];
@(posedge clk);
#1;data_in = testData6[4174];
@(posedge clk);
#1;data_in = testData6[4175];
@(posedge clk);
#1;data_in = testData6[4176];
@(posedge clk);
#1;data_in = testData6[4177];
@(posedge clk);
#1;data_in = testData6[4178];
@(posedge clk);
#1;data_in = testData6[4179];
@(posedge clk);
#1;data_in = testData6[4180];
@(posedge clk);
#1;data_in = testData6[4181];
@(posedge clk);
#1;data_in = testData6[4182];
@(posedge clk);
#1;data_in = testData6[4183];
@(posedge clk);
#1;data_in = testData6[4184];
@(posedge clk);
#1;data_in = testData6[4185];
@(posedge clk);
#1;data_in = testData6[4186];
@(posedge clk);
#1;data_in = testData6[4187];
@(posedge clk);
#1;data_in = testData6[4188];
@(posedge clk);
#1;data_in = testData6[4189];
@(posedge clk);
#1;data_in = testData6[4190];
@(posedge clk);
#1;data_in = testData6[4191];
@(posedge clk);
#1;data_in = testData6[4192];
@(posedge clk);
#1;data_in = testData6[4193];
@(posedge clk);
#1;data_in = testData6[4194];
@(posedge clk);
#1;data_in = testData6[4195];
@(posedge clk);
#1;data_in = testData6[4196];
@(posedge clk);
#1;data_in = testData6[4197];
@(posedge clk);
#1;data_in = testData6[4198];
@(posedge clk);
#1;data_in = testData6[4199];
@(posedge clk);
#1;data_in = testData6[4200];
@(posedge clk);
#1;data_in = testData6[4201];
@(posedge clk);
#1;data_in = testData6[4202];
@(posedge clk);
#1;data_in = testData6[4203];
@(posedge clk);
#1;data_in = testData6[4204];
@(posedge clk);
#1;data_in = testData6[4205];
@(posedge clk);
#1;data_in = testData6[4206];
@(posedge clk);
#1;data_in = testData6[4207];
@(posedge clk);
#1;data_in = testData6[4208];
@(posedge clk);
#1;data_in = testData6[4209];
@(posedge clk);
#1;data_in = testData6[4210];
@(posedge clk);
#1;data_in = testData6[4211];
@(posedge clk);
#1;data_in = testData6[4212];
@(posedge clk);
#1;data_in = testData6[4213];
@(posedge clk);
#1;data_in = testData6[4214];
@(posedge clk);
#1;data_in = testData6[4215];
@(posedge clk);
#1;data_in = testData6[4216];
@(posedge clk);
#1;data_in = testData6[4217];
@(posedge clk);
#1;data_in = testData6[4218];
@(posedge clk);
#1;data_in = testData6[4219];
@(posedge clk);
#1;data_in = testData6[4220];
@(posedge clk);
#1;data_in = testData6[4221];
@(posedge clk);
#1;data_in = testData6[4222];
@(posedge clk);
#1;data_in = testData6[4223];
@(posedge clk);
#1;data_in = testData6[4224];
@(posedge clk);
#1;data_in = testData6[4225];
@(posedge clk);
#1;data_in = testData6[4226];
@(posedge clk);
#1;data_in = testData6[4227];
@(posedge clk);
#1;data_in = testData6[4228];
@(posedge clk);
#1;data_in = testData6[4229];
@(posedge clk);
#1;data_in = testData6[4230];
@(posedge clk);
#1;data_in = testData6[4231];
@(posedge clk);
#1;data_in = testData6[4232];
@(posedge clk);
#1;data_in = testData6[4233];
@(posedge clk);
#1;data_in = testData6[4234];
@(posedge clk);
#1;data_in = testData6[4235];
@(posedge clk);
#1;data_in = testData6[4236];
@(posedge clk);
#1;data_in = testData6[4237];
@(posedge clk);
#1;data_in = testData6[4238];
@(posedge clk);
#1;data_in = testData6[4239];
@(posedge clk);
#1;data_in = testData6[4240];
@(posedge clk);
#1;data_in = testData6[4241];
@(posedge clk);
#1;data_in = testData6[4242];
@(posedge clk);
#1;data_in = testData6[4243];
@(posedge clk);
#1;data_in = testData6[4244];
@(posedge clk);
#1;data_in = testData6[4245];
@(posedge clk);
#1;data_in = testData6[4246];
@(posedge clk);
#1;data_in = testData6[4247];
@(posedge clk);
#1;data_in = testData6[4248];
@(posedge clk);
#1;data_in = testData6[4249];
@(posedge clk);
#1;data_in = testData6[4250];
@(posedge clk);
#1;data_in = testData6[4251];
@(posedge clk);
#1;data_in = testData6[4252];
@(posedge clk);
#1;data_in = testData6[4253];
@(posedge clk);
#1;data_in = testData6[4254];
@(posedge clk);
#1;data_in = testData6[4255];
@(posedge clk);
#1;data_in = testData6[4256];
@(posedge clk);
#1;data_in = testData6[4257];
@(posedge clk);
#1;data_in = testData6[4258];
@(posedge clk);
#1;data_in = testData6[4259];
@(posedge clk);
#1;data_in = testData6[4260];
@(posedge clk);
#1;data_in = testData6[4261];
@(posedge clk);
#1;data_in = testData6[4262];
@(posedge clk);
#1;data_in = testData6[4263];
@(posedge clk);
#1;data_in = testData6[4264];
@(posedge clk);
#1;data_in = testData6[4265];
@(posedge clk);
#1;data_in = testData6[4266];
@(posedge clk);
#1;data_in = testData6[4267];
@(posedge clk);
#1;data_in = testData6[4268];
@(posedge clk);
#1;data_in = testData6[4269];
@(posedge clk);
#1;data_in = testData6[4270];
@(posedge clk);
#1;data_in = testData6[4271];
@(posedge clk);
#1;data_in = testData6[4272];
@(posedge clk);
#1;data_in = testData6[4273];
@(posedge clk);
#1;data_in = testData6[4274];
@(posedge clk);
#1;data_in = testData6[4275];
@(posedge clk);
#1;data_in = testData6[4276];
@(posedge clk);
#1;data_in = testData6[4277];
@(posedge clk);
#1;data_in = testData6[4278];
@(posedge clk);
#1;data_in = testData6[4279];
@(posedge clk);
#1;data_in = testData6[4280];
@(posedge clk);
#1;data_in = testData6[4281];
@(posedge clk);
#1;data_in = testData6[4282];
@(posedge clk);
#1;data_in = testData6[4283];
@(posedge clk);
#1;data_in = testData6[4284];
@(posedge clk);
#1;data_in = testData6[4285];
@(posedge clk);
#1;data_in = testData6[4286];
@(posedge clk);
#1;data_in = testData6[4287];
@(posedge clk);
#1;data_in = testData6[4288];
@(posedge clk);
#1;data_in = testData6[4289];
@(posedge clk);
#1;data_in = testData6[4290];
@(posedge clk);
#1;data_in = testData6[4291];
@(posedge clk);
#1;data_in = testData6[4292];
@(posedge clk);
#1;data_in = testData6[4293];
@(posedge clk);
#1;data_in = testData6[4294];
@(posedge clk);
#1;data_in = testData6[4295];
@(posedge clk);
#1;data_in = testData6[4296];
@(posedge clk);
#1;data_in = testData6[4297];
@(posedge clk);
#1;data_in = testData6[4298];
@(posedge clk);
#1;data_in = testData6[4299];
@(posedge clk);
#1;data_in = testData6[4300];
@(posedge clk);
#1;data_in = testData6[4301];
@(posedge clk);
#1;data_in = testData6[4302];
@(posedge clk);
#1;data_in = testData6[4303];
@(posedge clk);
#1;data_in = testData6[4304];
@(posedge clk);
#1;data_in = testData6[4305];
@(posedge clk);
#1;data_in = testData6[4306];
@(posedge clk);
#1;data_in = testData6[4307];
@(posedge clk);
#1;data_in = testData6[4308];
@(posedge clk);
#1;data_in = testData6[4309];
@(posedge clk);
#1;data_in = testData6[4310];
@(posedge clk);
#1;data_in = testData6[4311];
@(posedge clk);
#1;data_in = testData6[4312];
@(posedge clk);
#1;data_in = testData6[4313];
@(posedge clk);
#1;data_in = testData6[4314];
@(posedge clk);
#1;data_in = testData6[4315];
@(posedge clk);
#1;data_in = testData6[4316];
@(posedge clk);
#1;data_in = testData6[4317];
@(posedge clk);
#1;data_in = testData6[4318];
@(posedge clk);
#1;data_in = testData6[4319];
@(posedge clk);
#1;data_in = testData6[4320];
@(posedge clk);
#1;data_in = testData6[4321];
@(posedge clk);
#1;data_in = testData6[4322];
@(posedge clk);
#1;data_in = testData6[4323];
@(posedge clk);
#1;data_in = testData6[4324];
@(posedge clk);
#1;data_in = testData6[4325];
@(posedge clk);
#1;data_in = testData6[4326];
@(posedge clk);
#1;data_in = testData6[4327];
@(posedge clk);
#1;data_in = testData6[4328];
@(posedge clk);
#1;data_in = testData6[4329];
@(posedge clk);
#1;data_in = testData6[4330];
@(posedge clk);
#1;data_in = testData6[4331];
@(posedge clk);
#1;data_in = testData6[4332];
@(posedge clk);
#1;data_in = testData6[4333];
@(posedge clk);
#1;data_in = testData6[4334];
@(posedge clk);
#1;data_in = testData6[4335];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[4336]; 
@(posedge clk);
#1;data_in = testData6[4337];
@(posedge clk);
#1;data_in = testData6[4338];
@(posedge clk);
#1;data_in = testData6[4339];
@(posedge clk);
#1;data_in = testData6[4340];
@(posedge clk);
#1;data_in = testData6[4341];
@(posedge clk);
#1;data_in = testData6[4342];
@(posedge clk);
#1;data_in = testData6[4343];
@(posedge clk);
#1;data_in = testData6[4344];
@(posedge clk);
#1;data_in = testData6[4345];
@(posedge clk);
#1;data_in = testData6[4346];
@(posedge clk);
#1;data_in = testData6[4347];
@(posedge clk);
#1;data_in = testData6[4348];
@(posedge clk);
#1;data_in = testData6[4349];
@(posedge clk);
#1;data_in = testData6[4350];
@(posedge clk);
#1;data_in = testData6[4351];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[4352];
@(posedge clk);
#1;data_in = testData6[4353];
@(posedge clk);
#1;data_in = testData6[4354];
@(posedge clk);
#1;data_in = testData6[4355];
@(posedge clk);
#1;data_in = testData6[4356];
@(posedge clk);
#1;data_in = testData6[4357];
@(posedge clk);
#1;data_in = testData6[4358];
@(posedge clk);
#1;data_in = testData6[4359];
@(posedge clk);
#1;data_in = testData6[4360];
@(posedge clk);
#1;data_in = testData6[4361];
@(posedge clk);
#1;data_in = testData6[4362];
@(posedge clk);
#1;data_in = testData6[4363];
@(posedge clk);
#1;data_in = testData6[4364];
@(posedge clk);
#1;data_in = testData6[4365];
@(posedge clk);
#1;data_in = testData6[4366];
@(posedge clk);
#1;data_in = testData6[4367];
@(posedge clk);
#1;data_in = testData6[4368];
@(posedge clk);
#1;data_in = testData6[4369];
@(posedge clk);
#1;data_in = testData6[4370];
@(posedge clk);
#1;data_in = testData6[4371];
@(posedge clk);
#1;data_in = testData6[4372];
@(posedge clk);
#1;data_in = testData6[4373];
@(posedge clk);
#1;data_in = testData6[4374];
@(posedge clk);
#1;data_in = testData6[4375];
@(posedge clk);
#1;data_in = testData6[4376];
@(posedge clk);
#1;data_in = testData6[4377];
@(posedge clk);
#1;data_in = testData6[4378];
@(posedge clk);
#1;data_in = testData6[4379];
@(posedge clk);
#1;data_in = testData6[4380];
@(posedge clk);
#1;data_in = testData6[4381];
@(posedge clk);
#1;data_in = testData6[4382];
@(posedge clk);
#1;data_in = testData6[4383];
@(posedge clk);
#1;data_in = testData6[4384];
@(posedge clk);
#1;data_in = testData6[4385];
@(posedge clk);
#1;data_in = testData6[4386];
@(posedge clk);
#1;data_in = testData6[4387];
@(posedge clk);
#1;data_in = testData6[4388];
@(posedge clk);
#1;data_in = testData6[4389];
@(posedge clk);
#1;data_in = testData6[4390];
@(posedge clk);
#1;data_in = testData6[4391];
@(posedge clk);
#1;data_in = testData6[4392];
@(posedge clk);
#1;data_in = testData6[4393];
@(posedge clk);
#1;data_in = testData6[4394];
@(posedge clk);
#1;data_in = testData6[4395];
@(posedge clk);
#1;data_in = testData6[4396];
@(posedge clk);
#1;data_in = testData6[4397];
@(posedge clk);
#1;data_in = testData6[4398];
@(posedge clk);
#1;data_in = testData6[4399];
@(posedge clk);
#1;data_in = testData6[4400];
@(posedge clk);
#1;data_in = testData6[4401];
@(posedge clk);
#1;data_in = testData6[4402];
@(posedge clk);
#1;data_in = testData6[4403];
@(posedge clk);
#1;data_in = testData6[4404];
@(posedge clk);
#1;data_in = testData6[4405];
@(posedge clk);
#1;data_in = testData6[4406];
@(posedge clk);
#1;data_in = testData6[4407];
@(posedge clk);
#1;data_in = testData6[4408];
@(posedge clk);
#1;data_in = testData6[4409];
@(posedge clk);
#1;data_in = testData6[4410];
@(posedge clk);
#1;data_in = testData6[4411];
@(posedge clk);
#1;data_in = testData6[4412];
@(posedge clk);
#1;data_in = testData6[4413];
@(posedge clk);
#1;data_in = testData6[4414];
@(posedge clk);
#1;data_in = testData6[4415];
@(posedge clk);
#1;data_in = testData6[4416];
@(posedge clk);
#1;data_in = testData6[4417];
@(posedge clk);
#1;data_in = testData6[4418];
@(posedge clk);
#1;data_in = testData6[4419];
@(posedge clk);
#1;data_in = testData6[4420];
@(posedge clk);
#1;data_in = testData6[4421];
@(posedge clk);
#1;data_in = testData6[4422];
@(posedge clk);
#1;data_in = testData6[4423];
@(posedge clk);
#1;data_in = testData6[4424];
@(posedge clk);
#1;data_in = testData6[4425];
@(posedge clk);
#1;data_in = testData6[4426];
@(posedge clk);
#1;data_in = testData6[4427];
@(posedge clk);
#1;data_in = testData6[4428];
@(posedge clk);
#1;data_in = testData6[4429];
@(posedge clk);
#1;data_in = testData6[4430];
@(posedge clk);
#1;data_in = testData6[4431];
@(posedge clk);
#1;data_in = testData6[4432];
@(posedge clk);
#1;data_in = testData6[4433];
@(posedge clk);
#1;data_in = testData6[4434];
@(posedge clk);
#1;data_in = testData6[4435];
@(posedge clk);
#1;data_in = testData6[4436];
@(posedge clk);
#1;data_in = testData6[4437];
@(posedge clk);
#1;data_in = testData6[4438];
@(posedge clk);
#1;data_in = testData6[4439];
@(posedge clk);
#1;data_in = testData6[4440];
@(posedge clk);
#1;data_in = testData6[4441];
@(posedge clk);
#1;data_in = testData6[4442];
@(posedge clk);
#1;data_in = testData6[4443];
@(posedge clk);
#1;data_in = testData6[4444];
@(posedge clk);
#1;data_in = testData6[4445];
@(posedge clk);
#1;data_in = testData6[4446];
@(posedge clk);
#1;data_in = testData6[4447];
@(posedge clk);
#1;data_in = testData6[4448];
@(posedge clk);
#1;data_in = testData6[4449];
@(posedge clk);
#1;data_in = testData6[4450];
@(posedge clk);
#1;data_in = testData6[4451];
@(posedge clk);
#1;data_in = testData6[4452];
@(posedge clk);
#1;data_in = testData6[4453];
@(posedge clk);
#1;data_in = testData6[4454];
@(posedge clk);
#1;data_in = testData6[4455];
@(posedge clk);
#1;data_in = testData6[4456];
@(posedge clk);
#1;data_in = testData6[4457];
@(posedge clk);
#1;data_in = testData6[4458];
@(posedge clk);
#1;data_in = testData6[4459];
@(posedge clk);
#1;data_in = testData6[4460];
@(posedge clk);
#1;data_in = testData6[4461];
@(posedge clk);
#1;data_in = testData6[4462];
@(posedge clk);
#1;data_in = testData6[4463];
@(posedge clk);
#1;data_in = testData6[4464];
@(posedge clk);
#1;data_in = testData6[4465];
@(posedge clk);
#1;data_in = testData6[4466];
@(posedge clk);
#1;data_in = testData6[4467];
@(posedge clk);
#1;data_in = testData6[4468];
@(posedge clk);
#1;data_in = testData6[4469];
@(posedge clk);
#1;data_in = testData6[4470];
@(posedge clk);
#1;data_in = testData6[4471];
@(posedge clk);
#1;data_in = testData6[4472];
@(posedge clk);
#1;data_in = testData6[4473];
@(posedge clk);
#1;data_in = testData6[4474];
@(posedge clk);
#1;data_in = testData6[4475];
@(posedge clk);
#1;data_in = testData6[4476];
@(posedge clk);
#1;data_in = testData6[4477];
@(posedge clk);
#1;data_in = testData6[4478];
@(posedge clk);
#1;data_in = testData6[4479];
@(posedge clk);
#1;data_in = testData6[4480];
@(posedge clk);
#1;data_in = testData6[4481];
@(posedge clk);
#1;data_in = testData6[4482];
@(posedge clk);
#1;data_in = testData6[4483];
@(posedge clk);
#1;data_in = testData6[4484];
@(posedge clk);
#1;data_in = testData6[4485];
@(posedge clk);
#1;data_in = testData6[4486];
@(posedge clk);
#1;data_in = testData6[4487];
@(posedge clk);
#1;data_in = testData6[4488];
@(posedge clk);
#1;data_in = testData6[4489];
@(posedge clk);
#1;data_in = testData6[4490];
@(posedge clk);
#1;data_in = testData6[4491];
@(posedge clk);
#1;data_in = testData6[4492];
@(posedge clk);
#1;data_in = testData6[4493];
@(posedge clk);
#1;data_in = testData6[4494];
@(posedge clk);
#1;data_in = testData6[4495];
@(posedge clk);
#1;data_in = testData6[4496];
@(posedge clk);
#1;data_in = testData6[4497];
@(posedge clk);
#1;data_in = testData6[4498];
@(posedge clk);
#1;data_in = testData6[4499];
@(posedge clk);
#1;data_in = testData6[4500];
@(posedge clk);
#1;data_in = testData6[4501];
@(posedge clk);
#1;data_in = testData6[4502];
@(posedge clk);
#1;data_in = testData6[4503];
@(posedge clk);
#1;data_in = testData6[4504];
@(posedge clk);
#1;data_in = testData6[4505];
@(posedge clk);
#1;data_in = testData6[4506];
@(posedge clk);
#1;data_in = testData6[4507];
@(posedge clk);
#1;data_in = testData6[4508];
@(posedge clk);
#1;data_in = testData6[4509];
@(posedge clk);
#1;data_in = testData6[4510];
@(posedge clk);
#1;data_in = testData6[4511];
@(posedge clk);
#1;data_in = testData6[4512];
@(posedge clk);
#1;data_in = testData6[4513];
@(posedge clk);
#1;data_in = testData6[4514];
@(posedge clk);
#1;data_in = testData6[4515];
@(posedge clk);
#1;data_in = testData6[4516];
@(posedge clk);
#1;data_in = testData6[4517];
@(posedge clk);
#1;data_in = testData6[4518];
@(posedge clk);
#1;data_in = testData6[4519];
@(posedge clk);
#1;data_in = testData6[4520];
@(posedge clk);
#1;data_in = testData6[4521];
@(posedge clk);
#1;data_in = testData6[4522];
@(posedge clk);
#1;data_in = testData6[4523];
@(posedge clk);
#1;data_in = testData6[4524];
@(posedge clk);
#1;data_in = testData6[4525];
@(posedge clk);
#1;data_in = testData6[4526];
@(posedge clk);
#1;data_in = testData6[4527];
@(posedge clk);
#1;data_in = testData6[4528];
@(posedge clk);
#1;data_in = testData6[4529];
@(posedge clk);
#1;data_in = testData6[4530];
@(posedge clk);
#1;data_in = testData6[4531];
@(posedge clk);
#1;data_in = testData6[4532];
@(posedge clk);
#1;data_in = testData6[4533];
@(posedge clk);
#1;data_in = testData6[4534];
@(posedge clk);
#1;data_in = testData6[4535];
@(posedge clk);
#1;data_in = testData6[4536];
@(posedge clk);
#1;data_in = testData6[4537];
@(posedge clk);
#1;data_in = testData6[4538];
@(posedge clk);
#1;data_in = testData6[4539];
@(posedge clk);
#1;data_in = testData6[4540];
@(posedge clk);
#1;data_in = testData6[4541];
@(posedge clk);
#1;data_in = testData6[4542];
@(posedge clk);
#1;data_in = testData6[4543];
@(posedge clk);
#1;data_in = testData6[4544];
@(posedge clk);
#1;data_in = testData6[4545];
@(posedge clk);
#1;data_in = testData6[4546];
@(posedge clk);
#1;data_in = testData6[4547];
@(posedge clk);
#1;data_in = testData6[4548];
@(posedge clk);
#1;data_in = testData6[4549];
@(posedge clk);
#1;data_in = testData6[4550];
@(posedge clk);
#1;data_in = testData6[4551];
@(posedge clk);
#1;data_in = testData6[4552];
@(posedge clk);
#1;data_in = testData6[4553];
@(posedge clk);
#1;data_in = testData6[4554];
@(posedge clk);
#1;data_in = testData6[4555];
@(posedge clk);
#1;data_in = testData6[4556];
@(posedge clk);
#1;data_in = testData6[4557];
@(posedge clk);
#1;data_in = testData6[4558];
@(posedge clk);
#1;data_in = testData6[4559];
@(posedge clk);
#1;data_in = testData6[4560];
@(posedge clk);
#1;data_in = testData6[4561];
@(posedge clk);
#1;data_in = testData6[4562];
@(posedge clk);
#1;data_in = testData6[4563];
@(posedge clk);
#1;data_in = testData6[4564];
@(posedge clk);
#1;data_in = testData6[4565];
@(posedge clk);
#1;data_in = testData6[4566];
@(posedge clk);
#1;data_in = testData6[4567];
@(posedge clk);
#1;data_in = testData6[4568];
@(posedge clk);
#1;data_in = testData6[4569];
@(posedge clk);
#1;data_in = testData6[4570];
@(posedge clk);
#1;data_in = testData6[4571];
@(posedge clk);
#1;data_in = testData6[4572];
@(posedge clk);
#1;data_in = testData6[4573];
@(posedge clk);
#1;data_in = testData6[4574];
@(posedge clk);
#1;data_in = testData6[4575];
@(posedge clk);
#1;data_in = testData6[4576];
@(posedge clk);
#1;data_in = testData6[4577];
@(posedge clk);
#1;data_in = testData6[4578];
@(posedge clk);
#1;data_in = testData6[4579];
@(posedge clk);
#1;data_in = testData6[4580];
@(posedge clk);
#1;data_in = testData6[4581];
@(posedge clk);
#1;data_in = testData6[4582];
@(posedge clk);
#1;data_in = testData6[4583];
@(posedge clk);
#1;data_in = testData6[4584];
@(posedge clk);
#1;data_in = testData6[4585];
@(posedge clk);
#1;data_in = testData6[4586];
@(posedge clk);
#1;data_in = testData6[4587];
@(posedge clk);
#1;data_in = testData6[4588];
@(posedge clk);
#1;data_in = testData6[4589];
@(posedge clk);
#1;data_in = testData6[4590];
@(posedge clk);
#1;data_in = testData6[4591];
@(posedge clk);
#1;data_in = testData6[4592];
@(posedge clk);
#1;data_in = testData6[4593];
@(posedge clk);
#1;data_in = testData6[4594];
@(posedge clk);
#1;data_in = testData6[4595];
@(posedge clk);
#1;data_in = testData6[4596];
@(posedge clk);
#1;data_in = testData6[4597];
@(posedge clk);
#1;data_in = testData6[4598];
@(posedge clk);
#1;data_in = testData6[4599];
@(posedge clk);
#1;data_in = testData6[4600];
@(posedge clk);
#1;data_in = testData6[4601];
@(posedge clk);
#1;data_in = testData6[4602];
@(posedge clk);
#1;data_in = testData6[4603];
@(posedge clk);
#1;data_in = testData6[4604];
@(posedge clk);
#1;data_in = testData6[4605];
@(posedge clk);
#1;data_in = testData6[4606];
@(posedge clk);
#1;data_in = testData6[4607];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[4608]; 
@(posedge clk);
#1;data_in = testData6[4609];
@(posedge clk);
#1;data_in = testData6[4610];
@(posedge clk);
#1;data_in = testData6[4611];
@(posedge clk);
#1;data_in = testData6[4612];
@(posedge clk);
#1;data_in = testData6[4613];
@(posedge clk);
#1;data_in = testData6[4614];
@(posedge clk);
#1;data_in = testData6[4615];
@(posedge clk);
#1;data_in = testData6[4616];
@(posedge clk);
#1;data_in = testData6[4617];
@(posedge clk);
#1;data_in = testData6[4618];
@(posedge clk);
#1;data_in = testData6[4619];
@(posedge clk);
#1;data_in = testData6[4620];
@(posedge clk);
#1;data_in = testData6[4621];
@(posedge clk);
#1;data_in = testData6[4622];
@(posedge clk);
#1;data_in = testData6[4623];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[4624];
@(posedge clk);
#1;data_in = testData6[4625];
@(posedge clk);
#1;data_in = testData6[4626];
@(posedge clk);
#1;data_in = testData6[4627];
@(posedge clk);
#1;data_in = testData6[4628];
@(posedge clk);
#1;data_in = testData6[4629];
@(posedge clk);
#1;data_in = testData6[4630];
@(posedge clk);
#1;data_in = testData6[4631];
@(posedge clk);
#1;data_in = testData6[4632];
@(posedge clk);
#1;data_in = testData6[4633];
@(posedge clk);
#1;data_in = testData6[4634];
@(posedge clk);
#1;data_in = testData6[4635];
@(posedge clk);
#1;data_in = testData6[4636];
@(posedge clk);
#1;data_in = testData6[4637];
@(posedge clk);
#1;data_in = testData6[4638];
@(posedge clk);
#1;data_in = testData6[4639];
@(posedge clk);
#1;data_in = testData6[4640];
@(posedge clk);
#1;data_in = testData6[4641];
@(posedge clk);
#1;data_in = testData6[4642];
@(posedge clk);
#1;data_in = testData6[4643];
@(posedge clk);
#1;data_in = testData6[4644];
@(posedge clk);
#1;data_in = testData6[4645];
@(posedge clk);
#1;data_in = testData6[4646];
@(posedge clk);
#1;data_in = testData6[4647];
@(posedge clk);
#1;data_in = testData6[4648];
@(posedge clk);
#1;data_in = testData6[4649];
@(posedge clk);
#1;data_in = testData6[4650];
@(posedge clk);
#1;data_in = testData6[4651];
@(posedge clk);
#1;data_in = testData6[4652];
@(posedge clk);
#1;data_in = testData6[4653];
@(posedge clk);
#1;data_in = testData6[4654];
@(posedge clk);
#1;data_in = testData6[4655];
@(posedge clk);
#1;data_in = testData6[4656];
@(posedge clk);
#1;data_in = testData6[4657];
@(posedge clk);
#1;data_in = testData6[4658];
@(posedge clk);
#1;data_in = testData6[4659];
@(posedge clk);
#1;data_in = testData6[4660];
@(posedge clk);
#1;data_in = testData6[4661];
@(posedge clk);
#1;data_in = testData6[4662];
@(posedge clk);
#1;data_in = testData6[4663];
@(posedge clk);
#1;data_in = testData6[4664];
@(posedge clk);
#1;data_in = testData6[4665];
@(posedge clk);
#1;data_in = testData6[4666];
@(posedge clk);
#1;data_in = testData6[4667];
@(posedge clk);
#1;data_in = testData6[4668];
@(posedge clk);
#1;data_in = testData6[4669];
@(posedge clk);
#1;data_in = testData6[4670];
@(posedge clk);
#1;data_in = testData6[4671];
@(posedge clk);
#1;data_in = testData6[4672];
@(posedge clk);
#1;data_in = testData6[4673];
@(posedge clk);
#1;data_in = testData6[4674];
@(posedge clk);
#1;data_in = testData6[4675];
@(posedge clk);
#1;data_in = testData6[4676];
@(posedge clk);
#1;data_in = testData6[4677];
@(posedge clk);
#1;data_in = testData6[4678];
@(posedge clk);
#1;data_in = testData6[4679];
@(posedge clk);
#1;data_in = testData6[4680];
@(posedge clk);
#1;data_in = testData6[4681];
@(posedge clk);
#1;data_in = testData6[4682];
@(posedge clk);
#1;data_in = testData6[4683];
@(posedge clk);
#1;data_in = testData6[4684];
@(posedge clk);
#1;data_in = testData6[4685];
@(posedge clk);
#1;data_in = testData6[4686];
@(posedge clk);
#1;data_in = testData6[4687];
@(posedge clk);
#1;data_in = testData6[4688];
@(posedge clk);
#1;data_in = testData6[4689];
@(posedge clk);
#1;data_in = testData6[4690];
@(posedge clk);
#1;data_in = testData6[4691];
@(posedge clk);
#1;data_in = testData6[4692];
@(posedge clk);
#1;data_in = testData6[4693];
@(posedge clk);
#1;data_in = testData6[4694];
@(posedge clk);
#1;data_in = testData6[4695];
@(posedge clk);
#1;data_in = testData6[4696];
@(posedge clk);
#1;data_in = testData6[4697];
@(posedge clk);
#1;data_in = testData6[4698];
@(posedge clk);
#1;data_in = testData6[4699];
@(posedge clk);
#1;data_in = testData6[4700];
@(posedge clk);
#1;data_in = testData6[4701];
@(posedge clk);
#1;data_in = testData6[4702];
@(posedge clk);
#1;data_in = testData6[4703];
@(posedge clk);
#1;data_in = testData6[4704];
@(posedge clk);
#1;data_in = testData6[4705];
@(posedge clk);
#1;data_in = testData6[4706];
@(posedge clk);
#1;data_in = testData6[4707];
@(posedge clk);
#1;data_in = testData6[4708];
@(posedge clk);
#1;data_in = testData6[4709];
@(posedge clk);
#1;data_in = testData6[4710];
@(posedge clk);
#1;data_in = testData6[4711];
@(posedge clk);
#1;data_in = testData6[4712];
@(posedge clk);
#1;data_in = testData6[4713];
@(posedge clk);
#1;data_in = testData6[4714];
@(posedge clk);
#1;data_in = testData6[4715];
@(posedge clk);
#1;data_in = testData6[4716];
@(posedge clk);
#1;data_in = testData6[4717];
@(posedge clk);
#1;data_in = testData6[4718];
@(posedge clk);
#1;data_in = testData6[4719];
@(posedge clk);
#1;data_in = testData6[4720];
@(posedge clk);
#1;data_in = testData6[4721];
@(posedge clk);
#1;data_in = testData6[4722];
@(posedge clk);
#1;data_in = testData6[4723];
@(posedge clk);
#1;data_in = testData6[4724];
@(posedge clk);
#1;data_in = testData6[4725];
@(posedge clk);
#1;data_in = testData6[4726];
@(posedge clk);
#1;data_in = testData6[4727];
@(posedge clk);
#1;data_in = testData6[4728];
@(posedge clk);
#1;data_in = testData6[4729];
@(posedge clk);
#1;data_in = testData6[4730];
@(posedge clk);
#1;data_in = testData6[4731];
@(posedge clk);
#1;data_in = testData6[4732];
@(posedge clk);
#1;data_in = testData6[4733];
@(posedge clk);
#1;data_in = testData6[4734];
@(posedge clk);
#1;data_in = testData6[4735];
@(posedge clk);
#1;data_in = testData6[4736];
@(posedge clk);
#1;data_in = testData6[4737];
@(posedge clk);
#1;data_in = testData6[4738];
@(posedge clk);
#1;data_in = testData6[4739];
@(posedge clk);
#1;data_in = testData6[4740];
@(posedge clk);
#1;data_in = testData6[4741];
@(posedge clk);
#1;data_in = testData6[4742];
@(posedge clk);
#1;data_in = testData6[4743];
@(posedge clk);
#1;data_in = testData6[4744];
@(posedge clk);
#1;data_in = testData6[4745];
@(posedge clk);
#1;data_in = testData6[4746];
@(posedge clk);
#1;data_in = testData6[4747];
@(posedge clk);
#1;data_in = testData6[4748];
@(posedge clk);
#1;data_in = testData6[4749];
@(posedge clk);
#1;data_in = testData6[4750];
@(posedge clk);
#1;data_in = testData6[4751];
@(posedge clk);
#1;data_in = testData6[4752];
@(posedge clk);
#1;data_in = testData6[4753];
@(posedge clk);
#1;data_in = testData6[4754];
@(posedge clk);
#1;data_in = testData6[4755];
@(posedge clk);
#1;data_in = testData6[4756];
@(posedge clk);
#1;data_in = testData6[4757];
@(posedge clk);
#1;data_in = testData6[4758];
@(posedge clk);
#1;data_in = testData6[4759];
@(posedge clk);
#1;data_in = testData6[4760];
@(posedge clk);
#1;data_in = testData6[4761];
@(posedge clk);
#1;data_in = testData6[4762];
@(posedge clk);
#1;data_in = testData6[4763];
@(posedge clk);
#1;data_in = testData6[4764];
@(posedge clk);
#1;data_in = testData6[4765];
@(posedge clk);
#1;data_in = testData6[4766];
@(posedge clk);
#1;data_in = testData6[4767];
@(posedge clk);
#1;data_in = testData6[4768];
@(posedge clk);
#1;data_in = testData6[4769];
@(posedge clk);
#1;data_in = testData6[4770];
@(posedge clk);
#1;data_in = testData6[4771];
@(posedge clk);
#1;data_in = testData6[4772];
@(posedge clk);
#1;data_in = testData6[4773];
@(posedge clk);
#1;data_in = testData6[4774];
@(posedge clk);
#1;data_in = testData6[4775];
@(posedge clk);
#1;data_in = testData6[4776];
@(posedge clk);
#1;data_in = testData6[4777];
@(posedge clk);
#1;data_in = testData6[4778];
@(posedge clk);
#1;data_in = testData6[4779];
@(posedge clk);
#1;data_in = testData6[4780];
@(posedge clk);
#1;data_in = testData6[4781];
@(posedge clk);
#1;data_in = testData6[4782];
@(posedge clk);
#1;data_in = testData6[4783];
@(posedge clk);
#1;data_in = testData6[4784];
@(posedge clk);
#1;data_in = testData6[4785];
@(posedge clk);
#1;data_in = testData6[4786];
@(posedge clk);
#1;data_in = testData6[4787];
@(posedge clk);
#1;data_in = testData6[4788];
@(posedge clk);
#1;data_in = testData6[4789];
@(posedge clk);
#1;data_in = testData6[4790];
@(posedge clk);
#1;data_in = testData6[4791];
@(posedge clk);
#1;data_in = testData6[4792];
@(posedge clk);
#1;data_in = testData6[4793];
@(posedge clk);
#1;data_in = testData6[4794];
@(posedge clk);
#1;data_in = testData6[4795];
@(posedge clk);
#1;data_in = testData6[4796];
@(posedge clk);
#1;data_in = testData6[4797];
@(posedge clk);
#1;data_in = testData6[4798];
@(posedge clk);
#1;data_in = testData6[4799];
@(posedge clk);
#1;data_in = testData6[4800];
@(posedge clk);
#1;data_in = testData6[4801];
@(posedge clk);
#1;data_in = testData6[4802];
@(posedge clk);
#1;data_in = testData6[4803];
@(posedge clk);
#1;data_in = testData6[4804];
@(posedge clk);
#1;data_in = testData6[4805];
@(posedge clk);
#1;data_in = testData6[4806];
@(posedge clk);
#1;data_in = testData6[4807];
@(posedge clk);
#1;data_in = testData6[4808];
@(posedge clk);
#1;data_in = testData6[4809];
@(posedge clk);
#1;data_in = testData6[4810];
@(posedge clk);
#1;data_in = testData6[4811];
@(posedge clk);
#1;data_in = testData6[4812];
@(posedge clk);
#1;data_in = testData6[4813];
@(posedge clk);
#1;data_in = testData6[4814];
@(posedge clk);
#1;data_in = testData6[4815];
@(posedge clk);
#1;data_in = testData6[4816];
@(posedge clk);
#1;data_in = testData6[4817];
@(posedge clk);
#1;data_in = testData6[4818];
@(posedge clk);
#1;data_in = testData6[4819];
@(posedge clk);
#1;data_in = testData6[4820];
@(posedge clk);
#1;data_in = testData6[4821];
@(posedge clk);
#1;data_in = testData6[4822];
@(posedge clk);
#1;data_in = testData6[4823];
@(posedge clk);
#1;data_in = testData6[4824];
@(posedge clk);
#1;data_in = testData6[4825];
@(posedge clk);
#1;data_in = testData6[4826];
@(posedge clk);
#1;data_in = testData6[4827];
@(posedge clk);
#1;data_in = testData6[4828];
@(posedge clk);
#1;data_in = testData6[4829];
@(posedge clk);
#1;data_in = testData6[4830];
@(posedge clk);
#1;data_in = testData6[4831];
@(posedge clk);
#1;data_in = testData6[4832];
@(posedge clk);
#1;data_in = testData6[4833];
@(posedge clk);
#1;data_in = testData6[4834];
@(posedge clk);
#1;data_in = testData6[4835];
@(posedge clk);
#1;data_in = testData6[4836];
@(posedge clk);
#1;data_in = testData6[4837];
@(posedge clk);
#1;data_in = testData6[4838];
@(posedge clk);
#1;data_in = testData6[4839];
@(posedge clk);
#1;data_in = testData6[4840];
@(posedge clk);
#1;data_in = testData6[4841];
@(posedge clk);
#1;data_in = testData6[4842];
@(posedge clk);
#1;data_in = testData6[4843];
@(posedge clk);
#1;data_in = testData6[4844];
@(posedge clk);
#1;data_in = testData6[4845];
@(posedge clk);
#1;data_in = testData6[4846];
@(posedge clk);
#1;data_in = testData6[4847];
@(posedge clk);
#1;data_in = testData6[4848];
@(posedge clk);
#1;data_in = testData6[4849];
@(posedge clk);
#1;data_in = testData6[4850];
@(posedge clk);
#1;data_in = testData6[4851];
@(posedge clk);
#1;data_in = testData6[4852];
@(posedge clk);
#1;data_in = testData6[4853];
@(posedge clk);
#1;data_in = testData6[4854];
@(posedge clk);
#1;data_in = testData6[4855];
@(posedge clk);
#1;data_in = testData6[4856];
@(posedge clk);
#1;data_in = testData6[4857];
@(posedge clk);
#1;data_in = testData6[4858];
@(posedge clk);
#1;data_in = testData6[4859];
@(posedge clk);
#1;data_in = testData6[4860];
@(posedge clk);
#1;data_in = testData6[4861];
@(posedge clk);
#1;data_in = testData6[4862];
@(posedge clk);
#1;data_in = testData6[4863];
@(posedge clk);
#1;data_in = testData6[4864];
@(posedge clk);
#1;data_in = testData6[4865];
@(posedge clk);
#1;data_in = testData6[4866];
@(posedge clk);
#1;data_in = testData6[4867];
@(posedge clk);
#1;data_in = testData6[4868];
@(posedge clk);
#1;data_in = testData6[4869];
@(posedge clk);
#1;data_in = testData6[4870];
@(posedge clk);
#1;data_in = testData6[4871];
@(posedge clk);
#1;data_in = testData6[4872];
@(posedge clk);
#1;data_in = testData6[4873];
@(posedge clk);
#1;data_in = testData6[4874];
@(posedge clk);
#1;data_in = testData6[4875];
@(posedge clk);
#1;data_in = testData6[4876];
@(posedge clk);
#1;data_in = testData6[4877];
@(posedge clk);
#1;data_in = testData6[4878];
@(posedge clk);
#1;data_in = testData6[4879];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[4880]; 
@(posedge clk);
#1;data_in = testData6[4881];
@(posedge clk);
#1;data_in = testData6[4882];
@(posedge clk);
#1;data_in = testData6[4883];
@(posedge clk);
#1;data_in = testData6[4884];
@(posedge clk);
#1;data_in = testData6[4885];
@(posedge clk);
#1;data_in = testData6[4886];
@(posedge clk);
#1;data_in = testData6[4887];
@(posedge clk);
#1;data_in = testData6[4888];
@(posedge clk);
#1;data_in = testData6[4889];
@(posedge clk);
#1;data_in = testData6[4890];
@(posedge clk);
#1;data_in = testData6[4891];
@(posedge clk);
#1;data_in = testData6[4892];
@(posedge clk);
#1;data_in = testData6[4893];
@(posedge clk);
#1;data_in = testData6[4894];
@(posedge clk);
#1;data_in = testData6[4895];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[4896];
@(posedge clk);
#1;data_in = testData6[4897];
@(posedge clk);
#1;data_in = testData6[4898];
@(posedge clk);
#1;data_in = testData6[4899];
@(posedge clk);
#1;data_in = testData6[4900];
@(posedge clk);
#1;data_in = testData6[4901];
@(posedge clk);
#1;data_in = testData6[4902];
@(posedge clk);
#1;data_in = testData6[4903];
@(posedge clk);
#1;data_in = testData6[4904];
@(posedge clk);
#1;data_in = testData6[4905];
@(posedge clk);
#1;data_in = testData6[4906];
@(posedge clk);
#1;data_in = testData6[4907];
@(posedge clk);
#1;data_in = testData6[4908];
@(posedge clk);
#1;data_in = testData6[4909];
@(posedge clk);
#1;data_in = testData6[4910];
@(posedge clk);
#1;data_in = testData6[4911];
@(posedge clk);
#1;data_in = testData6[4912];
@(posedge clk);
#1;data_in = testData6[4913];
@(posedge clk);
#1;data_in = testData6[4914];
@(posedge clk);
#1;data_in = testData6[4915];
@(posedge clk);
#1;data_in = testData6[4916];
@(posedge clk);
#1;data_in = testData6[4917];
@(posedge clk);
#1;data_in = testData6[4918];
@(posedge clk);
#1;data_in = testData6[4919];
@(posedge clk);
#1;data_in = testData6[4920];
@(posedge clk);
#1;data_in = testData6[4921];
@(posedge clk);
#1;data_in = testData6[4922];
@(posedge clk);
#1;data_in = testData6[4923];
@(posedge clk);
#1;data_in = testData6[4924];
@(posedge clk);
#1;data_in = testData6[4925];
@(posedge clk);
#1;data_in = testData6[4926];
@(posedge clk);
#1;data_in = testData6[4927];
@(posedge clk);
#1;data_in = testData6[4928];
@(posedge clk);
#1;data_in = testData6[4929];
@(posedge clk);
#1;data_in = testData6[4930];
@(posedge clk);
#1;data_in = testData6[4931];
@(posedge clk);
#1;data_in = testData6[4932];
@(posedge clk);
#1;data_in = testData6[4933];
@(posedge clk);
#1;data_in = testData6[4934];
@(posedge clk);
#1;data_in = testData6[4935];
@(posedge clk);
#1;data_in = testData6[4936];
@(posedge clk);
#1;data_in = testData6[4937];
@(posedge clk);
#1;data_in = testData6[4938];
@(posedge clk);
#1;data_in = testData6[4939];
@(posedge clk);
#1;data_in = testData6[4940];
@(posedge clk);
#1;data_in = testData6[4941];
@(posedge clk);
#1;data_in = testData6[4942];
@(posedge clk);
#1;data_in = testData6[4943];
@(posedge clk);
#1;data_in = testData6[4944];
@(posedge clk);
#1;data_in = testData6[4945];
@(posedge clk);
#1;data_in = testData6[4946];
@(posedge clk);
#1;data_in = testData6[4947];
@(posedge clk);
#1;data_in = testData6[4948];
@(posedge clk);
#1;data_in = testData6[4949];
@(posedge clk);
#1;data_in = testData6[4950];
@(posedge clk);
#1;data_in = testData6[4951];
@(posedge clk);
#1;data_in = testData6[4952];
@(posedge clk);
#1;data_in = testData6[4953];
@(posedge clk);
#1;data_in = testData6[4954];
@(posedge clk);
#1;data_in = testData6[4955];
@(posedge clk);
#1;data_in = testData6[4956];
@(posedge clk);
#1;data_in = testData6[4957];
@(posedge clk);
#1;data_in = testData6[4958];
@(posedge clk);
#1;data_in = testData6[4959];
@(posedge clk);
#1;data_in = testData6[4960];
@(posedge clk);
#1;data_in = testData6[4961];
@(posedge clk);
#1;data_in = testData6[4962];
@(posedge clk);
#1;data_in = testData6[4963];
@(posedge clk);
#1;data_in = testData6[4964];
@(posedge clk);
#1;data_in = testData6[4965];
@(posedge clk);
#1;data_in = testData6[4966];
@(posedge clk);
#1;data_in = testData6[4967];
@(posedge clk);
#1;data_in = testData6[4968];
@(posedge clk);
#1;data_in = testData6[4969];
@(posedge clk);
#1;data_in = testData6[4970];
@(posedge clk);
#1;data_in = testData6[4971];
@(posedge clk);
#1;data_in = testData6[4972];
@(posedge clk);
#1;data_in = testData6[4973];
@(posedge clk);
#1;data_in = testData6[4974];
@(posedge clk);
#1;data_in = testData6[4975];
@(posedge clk);
#1;data_in = testData6[4976];
@(posedge clk);
#1;data_in = testData6[4977];
@(posedge clk);
#1;data_in = testData6[4978];
@(posedge clk);
#1;data_in = testData6[4979];
@(posedge clk);
#1;data_in = testData6[4980];
@(posedge clk);
#1;data_in = testData6[4981];
@(posedge clk);
#1;data_in = testData6[4982];
@(posedge clk);
#1;data_in = testData6[4983];
@(posedge clk);
#1;data_in = testData6[4984];
@(posedge clk);
#1;data_in = testData6[4985];
@(posedge clk);
#1;data_in = testData6[4986];
@(posedge clk);
#1;data_in = testData6[4987];
@(posedge clk);
#1;data_in = testData6[4988];
@(posedge clk);
#1;data_in = testData6[4989];
@(posedge clk);
#1;data_in = testData6[4990];
@(posedge clk);
#1;data_in = testData6[4991];
@(posedge clk);
#1;data_in = testData6[4992];
@(posedge clk);
#1;data_in = testData6[4993];
@(posedge clk);
#1;data_in = testData6[4994];
@(posedge clk);
#1;data_in = testData6[4995];
@(posedge clk);
#1;data_in = testData6[4996];
@(posedge clk);
#1;data_in = testData6[4997];
@(posedge clk);
#1;data_in = testData6[4998];
@(posedge clk);
#1;data_in = testData6[4999];
@(posedge clk);
#1;data_in = testData6[5000];
@(posedge clk);
#1;data_in = testData6[5001];
@(posedge clk);
#1;data_in = testData6[5002];
@(posedge clk);
#1;data_in = testData6[5003];
@(posedge clk);
#1;data_in = testData6[5004];
@(posedge clk);
#1;data_in = testData6[5005];
@(posedge clk);
#1;data_in = testData6[5006];
@(posedge clk);
#1;data_in = testData6[5007];
@(posedge clk);
#1;data_in = testData6[5008];
@(posedge clk);
#1;data_in = testData6[5009];
@(posedge clk);
#1;data_in = testData6[5010];
@(posedge clk);
#1;data_in = testData6[5011];
@(posedge clk);
#1;data_in = testData6[5012];
@(posedge clk);
#1;data_in = testData6[5013];
@(posedge clk);
#1;data_in = testData6[5014];
@(posedge clk);
#1;data_in = testData6[5015];
@(posedge clk);
#1;data_in = testData6[5016];
@(posedge clk);
#1;data_in = testData6[5017];
@(posedge clk);
#1;data_in = testData6[5018];
@(posedge clk);
#1;data_in = testData6[5019];
@(posedge clk);
#1;data_in = testData6[5020];
@(posedge clk);
#1;data_in = testData6[5021];
@(posedge clk);
#1;data_in = testData6[5022];
@(posedge clk);
#1;data_in = testData6[5023];
@(posedge clk);
#1;data_in = testData6[5024];
@(posedge clk);
#1;data_in = testData6[5025];
@(posedge clk);
#1;data_in = testData6[5026];
@(posedge clk);
#1;data_in = testData6[5027];
@(posedge clk);
#1;data_in = testData6[5028];
@(posedge clk);
#1;data_in = testData6[5029];
@(posedge clk);
#1;data_in = testData6[5030];
@(posedge clk);
#1;data_in = testData6[5031];
@(posedge clk);
#1;data_in = testData6[5032];
@(posedge clk);
#1;data_in = testData6[5033];
@(posedge clk);
#1;data_in = testData6[5034];
@(posedge clk);
#1;data_in = testData6[5035];
@(posedge clk);
#1;data_in = testData6[5036];
@(posedge clk);
#1;data_in = testData6[5037];
@(posedge clk);
#1;data_in = testData6[5038];
@(posedge clk);
#1;data_in = testData6[5039];
@(posedge clk);
#1;data_in = testData6[5040];
@(posedge clk);
#1;data_in = testData6[5041];
@(posedge clk);
#1;data_in = testData6[5042];
@(posedge clk);
#1;data_in = testData6[5043];
@(posedge clk);
#1;data_in = testData6[5044];
@(posedge clk);
#1;data_in = testData6[5045];
@(posedge clk);
#1;data_in = testData6[5046];
@(posedge clk);
#1;data_in = testData6[5047];
@(posedge clk);
#1;data_in = testData6[5048];
@(posedge clk);
#1;data_in = testData6[5049];
@(posedge clk);
#1;data_in = testData6[5050];
@(posedge clk);
#1;data_in = testData6[5051];
@(posedge clk);
#1;data_in = testData6[5052];
@(posedge clk);
#1;data_in = testData6[5053];
@(posedge clk);
#1;data_in = testData6[5054];
@(posedge clk);
#1;data_in = testData6[5055];
@(posedge clk);
#1;data_in = testData6[5056];
@(posedge clk);
#1;data_in = testData6[5057];
@(posedge clk);
#1;data_in = testData6[5058];
@(posedge clk);
#1;data_in = testData6[5059];
@(posedge clk);
#1;data_in = testData6[5060];
@(posedge clk);
#1;data_in = testData6[5061];
@(posedge clk);
#1;data_in = testData6[5062];
@(posedge clk);
#1;data_in = testData6[5063];
@(posedge clk);
#1;data_in = testData6[5064];
@(posedge clk);
#1;data_in = testData6[5065];
@(posedge clk);
#1;data_in = testData6[5066];
@(posedge clk);
#1;data_in = testData6[5067];
@(posedge clk);
#1;data_in = testData6[5068];
@(posedge clk);
#1;data_in = testData6[5069];
@(posedge clk);
#1;data_in = testData6[5070];
@(posedge clk);
#1;data_in = testData6[5071];
@(posedge clk);
#1;data_in = testData6[5072];
@(posedge clk);
#1;data_in = testData6[5073];
@(posedge clk);
#1;data_in = testData6[5074];
@(posedge clk);
#1;data_in = testData6[5075];
@(posedge clk);
#1;data_in = testData6[5076];
@(posedge clk);
#1;data_in = testData6[5077];
@(posedge clk);
#1;data_in = testData6[5078];
@(posedge clk);
#1;data_in = testData6[5079];
@(posedge clk);
#1;data_in = testData6[5080];
@(posedge clk);
#1;data_in = testData6[5081];
@(posedge clk);
#1;data_in = testData6[5082];
@(posedge clk);
#1;data_in = testData6[5083];
@(posedge clk);
#1;data_in = testData6[5084];
@(posedge clk);
#1;data_in = testData6[5085];
@(posedge clk);
#1;data_in = testData6[5086];
@(posedge clk);
#1;data_in = testData6[5087];
@(posedge clk);
#1;data_in = testData6[5088];
@(posedge clk);
#1;data_in = testData6[5089];
@(posedge clk);
#1;data_in = testData6[5090];
@(posedge clk);
#1;data_in = testData6[5091];
@(posedge clk);
#1;data_in = testData6[5092];
@(posedge clk);
#1;data_in = testData6[5093];
@(posedge clk);
#1;data_in = testData6[5094];
@(posedge clk);
#1;data_in = testData6[5095];
@(posedge clk);
#1;data_in = testData6[5096];
@(posedge clk);
#1;data_in = testData6[5097];
@(posedge clk);
#1;data_in = testData6[5098];
@(posedge clk);
#1;data_in = testData6[5099];
@(posedge clk);
#1;data_in = testData6[5100];
@(posedge clk);
#1;data_in = testData6[5101];
@(posedge clk);
#1;data_in = testData6[5102];
@(posedge clk);
#1;data_in = testData6[5103];
@(posedge clk);
#1;data_in = testData6[5104];
@(posedge clk);
#1;data_in = testData6[5105];
@(posedge clk);
#1;data_in = testData6[5106];
@(posedge clk);
#1;data_in = testData6[5107];
@(posedge clk);
#1;data_in = testData6[5108];
@(posedge clk);
#1;data_in = testData6[5109];
@(posedge clk);
#1;data_in = testData6[5110];
@(posedge clk);
#1;data_in = testData6[5111];
@(posedge clk);
#1;data_in = testData6[5112];
@(posedge clk);
#1;data_in = testData6[5113];
@(posedge clk);
#1;data_in = testData6[5114];
@(posedge clk);
#1;data_in = testData6[5115];
@(posedge clk);
#1;data_in = testData6[5116];
@(posedge clk);
#1;data_in = testData6[5117];
@(posedge clk);
#1;data_in = testData6[5118];
@(posedge clk);
#1;data_in = testData6[5119];
@(posedge clk);
#1;data_in = testData6[5120];
@(posedge clk);
#1;data_in = testData6[5121];
@(posedge clk);
#1;data_in = testData6[5122];
@(posedge clk);
#1;data_in = testData6[5123];
@(posedge clk);
#1;data_in = testData6[5124];
@(posedge clk);
#1;data_in = testData6[5125];
@(posedge clk);
#1;data_in = testData6[5126];
@(posedge clk);
#1;data_in = testData6[5127];
@(posedge clk);
#1;data_in = testData6[5128];
@(posedge clk);
#1;data_in = testData6[5129];
@(posedge clk);
#1;data_in = testData6[5130];
@(posedge clk);
#1;data_in = testData6[5131];
@(posedge clk);
#1;data_in = testData6[5132];
@(posedge clk);
#1;data_in = testData6[5133];
@(posedge clk);
#1;data_in = testData6[5134];
@(posedge clk);
#1;data_in = testData6[5135];
@(posedge clk);
#1;data_in = testData6[5136];
@(posedge clk);
#1;data_in = testData6[5137];
@(posedge clk);
#1;data_in = testData6[5138];
@(posedge clk);
#1;data_in = testData6[5139];
@(posedge clk);
#1;data_in = testData6[5140];
@(posedge clk);
#1;data_in = testData6[5141];
@(posedge clk);
#1;data_in = testData6[5142];
@(posedge clk);
#1;data_in = testData6[5143];
@(posedge clk);
#1;data_in = testData6[5144];
@(posedge clk);
#1;data_in = testData6[5145];
@(posedge clk);
#1;data_in = testData6[5146];
@(posedge clk);
#1;data_in = testData6[5147];
@(posedge clk);
#1;data_in = testData6[5148];
@(posedge clk);
#1;data_in = testData6[5149];
@(posedge clk);
#1;data_in = testData6[5150];
@(posedge clk);
#1;data_in = testData6[5151];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[5152]; 
@(posedge clk);
#1;data_in = testData6[5153];
@(posedge clk);
#1;data_in = testData6[5154];
@(posedge clk);
#1;data_in = testData6[5155];
@(posedge clk);
#1;data_in = testData6[5156];
@(posedge clk);
#1;data_in = testData6[5157];
@(posedge clk);
#1;data_in = testData6[5158];
@(posedge clk);
#1;data_in = testData6[5159];
@(posedge clk);
#1;data_in = testData6[5160];
@(posedge clk);
#1;data_in = testData6[5161];
@(posedge clk);
#1;data_in = testData6[5162];
@(posedge clk);
#1;data_in = testData6[5163];
@(posedge clk);
#1;data_in = testData6[5164];
@(posedge clk);
#1;data_in = testData6[5165];
@(posedge clk);
#1;data_in = testData6[5166];
@(posedge clk);
#1;data_in = testData6[5167];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[5168];
@(posedge clk);
#1;data_in = testData6[5169];
@(posedge clk);
#1;data_in = testData6[5170];
@(posedge clk);
#1;data_in = testData6[5171];
@(posedge clk);
#1;data_in = testData6[5172];
@(posedge clk);
#1;data_in = testData6[5173];
@(posedge clk);
#1;data_in = testData6[5174];
@(posedge clk);
#1;data_in = testData6[5175];
@(posedge clk);
#1;data_in = testData6[5176];
@(posedge clk);
#1;data_in = testData6[5177];
@(posedge clk);
#1;data_in = testData6[5178];
@(posedge clk);
#1;data_in = testData6[5179];
@(posedge clk);
#1;data_in = testData6[5180];
@(posedge clk);
#1;data_in = testData6[5181];
@(posedge clk);
#1;data_in = testData6[5182];
@(posedge clk);
#1;data_in = testData6[5183];
@(posedge clk);
#1;data_in = testData6[5184];
@(posedge clk);
#1;data_in = testData6[5185];
@(posedge clk);
#1;data_in = testData6[5186];
@(posedge clk);
#1;data_in = testData6[5187];
@(posedge clk);
#1;data_in = testData6[5188];
@(posedge clk);
#1;data_in = testData6[5189];
@(posedge clk);
#1;data_in = testData6[5190];
@(posedge clk);
#1;data_in = testData6[5191];
@(posedge clk);
#1;data_in = testData6[5192];
@(posedge clk);
#1;data_in = testData6[5193];
@(posedge clk);
#1;data_in = testData6[5194];
@(posedge clk);
#1;data_in = testData6[5195];
@(posedge clk);
#1;data_in = testData6[5196];
@(posedge clk);
#1;data_in = testData6[5197];
@(posedge clk);
#1;data_in = testData6[5198];
@(posedge clk);
#1;data_in = testData6[5199];
@(posedge clk);
#1;data_in = testData6[5200];
@(posedge clk);
#1;data_in = testData6[5201];
@(posedge clk);
#1;data_in = testData6[5202];
@(posedge clk);
#1;data_in = testData6[5203];
@(posedge clk);
#1;data_in = testData6[5204];
@(posedge clk);
#1;data_in = testData6[5205];
@(posedge clk);
#1;data_in = testData6[5206];
@(posedge clk);
#1;data_in = testData6[5207];
@(posedge clk);
#1;data_in = testData6[5208];
@(posedge clk);
#1;data_in = testData6[5209];
@(posedge clk);
#1;data_in = testData6[5210];
@(posedge clk);
#1;data_in = testData6[5211];
@(posedge clk);
#1;data_in = testData6[5212];
@(posedge clk);
#1;data_in = testData6[5213];
@(posedge clk);
#1;data_in = testData6[5214];
@(posedge clk);
#1;data_in = testData6[5215];
@(posedge clk);
#1;data_in = testData6[5216];
@(posedge clk);
#1;data_in = testData6[5217];
@(posedge clk);
#1;data_in = testData6[5218];
@(posedge clk);
#1;data_in = testData6[5219];
@(posedge clk);
#1;data_in = testData6[5220];
@(posedge clk);
#1;data_in = testData6[5221];
@(posedge clk);
#1;data_in = testData6[5222];
@(posedge clk);
#1;data_in = testData6[5223];
@(posedge clk);
#1;data_in = testData6[5224];
@(posedge clk);
#1;data_in = testData6[5225];
@(posedge clk);
#1;data_in = testData6[5226];
@(posedge clk);
#1;data_in = testData6[5227];
@(posedge clk);
#1;data_in = testData6[5228];
@(posedge clk);
#1;data_in = testData6[5229];
@(posedge clk);
#1;data_in = testData6[5230];
@(posedge clk);
#1;data_in = testData6[5231];
@(posedge clk);
#1;data_in = testData6[5232];
@(posedge clk);
#1;data_in = testData6[5233];
@(posedge clk);
#1;data_in = testData6[5234];
@(posedge clk);
#1;data_in = testData6[5235];
@(posedge clk);
#1;data_in = testData6[5236];
@(posedge clk);
#1;data_in = testData6[5237];
@(posedge clk);
#1;data_in = testData6[5238];
@(posedge clk);
#1;data_in = testData6[5239];
@(posedge clk);
#1;data_in = testData6[5240];
@(posedge clk);
#1;data_in = testData6[5241];
@(posedge clk);
#1;data_in = testData6[5242];
@(posedge clk);
#1;data_in = testData6[5243];
@(posedge clk);
#1;data_in = testData6[5244];
@(posedge clk);
#1;data_in = testData6[5245];
@(posedge clk);
#1;data_in = testData6[5246];
@(posedge clk);
#1;data_in = testData6[5247];
@(posedge clk);
#1;data_in = testData6[5248];
@(posedge clk);
#1;data_in = testData6[5249];
@(posedge clk);
#1;data_in = testData6[5250];
@(posedge clk);
#1;data_in = testData6[5251];
@(posedge clk);
#1;data_in = testData6[5252];
@(posedge clk);
#1;data_in = testData6[5253];
@(posedge clk);
#1;data_in = testData6[5254];
@(posedge clk);
#1;data_in = testData6[5255];
@(posedge clk);
#1;data_in = testData6[5256];
@(posedge clk);
#1;data_in = testData6[5257];
@(posedge clk);
#1;data_in = testData6[5258];
@(posedge clk);
#1;data_in = testData6[5259];
@(posedge clk);
#1;data_in = testData6[5260];
@(posedge clk);
#1;data_in = testData6[5261];
@(posedge clk);
#1;data_in = testData6[5262];
@(posedge clk);
#1;data_in = testData6[5263];
@(posedge clk);
#1;data_in = testData6[5264];
@(posedge clk);
#1;data_in = testData6[5265];
@(posedge clk);
#1;data_in = testData6[5266];
@(posedge clk);
#1;data_in = testData6[5267];
@(posedge clk);
#1;data_in = testData6[5268];
@(posedge clk);
#1;data_in = testData6[5269];
@(posedge clk);
#1;data_in = testData6[5270];
@(posedge clk);
#1;data_in = testData6[5271];
@(posedge clk);
#1;data_in = testData6[5272];
@(posedge clk);
#1;data_in = testData6[5273];
@(posedge clk);
#1;data_in = testData6[5274];
@(posedge clk);
#1;data_in = testData6[5275];
@(posedge clk);
#1;data_in = testData6[5276];
@(posedge clk);
#1;data_in = testData6[5277];
@(posedge clk);
#1;data_in = testData6[5278];
@(posedge clk);
#1;data_in = testData6[5279];
@(posedge clk);
#1;data_in = testData6[5280];
@(posedge clk);
#1;data_in = testData6[5281];
@(posedge clk);
#1;data_in = testData6[5282];
@(posedge clk);
#1;data_in = testData6[5283];
@(posedge clk);
#1;data_in = testData6[5284];
@(posedge clk);
#1;data_in = testData6[5285];
@(posedge clk);
#1;data_in = testData6[5286];
@(posedge clk);
#1;data_in = testData6[5287];
@(posedge clk);
#1;data_in = testData6[5288];
@(posedge clk);
#1;data_in = testData6[5289];
@(posedge clk);
#1;data_in = testData6[5290];
@(posedge clk);
#1;data_in = testData6[5291];
@(posedge clk);
#1;data_in = testData6[5292];
@(posedge clk);
#1;data_in = testData6[5293];
@(posedge clk);
#1;data_in = testData6[5294];
@(posedge clk);
#1;data_in = testData6[5295];
@(posedge clk);
#1;data_in = testData6[5296];
@(posedge clk);
#1;data_in = testData6[5297];
@(posedge clk);
#1;data_in = testData6[5298];
@(posedge clk);
#1;data_in = testData6[5299];
@(posedge clk);
#1;data_in = testData6[5300];
@(posedge clk);
#1;data_in = testData6[5301];
@(posedge clk);
#1;data_in = testData6[5302];
@(posedge clk);
#1;data_in = testData6[5303];
@(posedge clk);
#1;data_in = testData6[5304];
@(posedge clk);
#1;data_in = testData6[5305];
@(posedge clk);
#1;data_in = testData6[5306];
@(posedge clk);
#1;data_in = testData6[5307];
@(posedge clk);
#1;data_in = testData6[5308];
@(posedge clk);
#1;data_in = testData6[5309];
@(posedge clk);
#1;data_in = testData6[5310];
@(posedge clk);
#1;data_in = testData6[5311];
@(posedge clk);
#1;data_in = testData6[5312];
@(posedge clk);
#1;data_in = testData6[5313];
@(posedge clk);
#1;data_in = testData6[5314];
@(posedge clk);
#1;data_in = testData6[5315];
@(posedge clk);
#1;data_in = testData6[5316];
@(posedge clk);
#1;data_in = testData6[5317];
@(posedge clk);
#1;data_in = testData6[5318];
@(posedge clk);
#1;data_in = testData6[5319];
@(posedge clk);
#1;data_in = testData6[5320];
@(posedge clk);
#1;data_in = testData6[5321];
@(posedge clk);
#1;data_in = testData6[5322];
@(posedge clk);
#1;data_in = testData6[5323];
@(posedge clk);
#1;data_in = testData6[5324];
@(posedge clk);
#1;data_in = testData6[5325];
@(posedge clk);
#1;data_in = testData6[5326];
@(posedge clk);
#1;data_in = testData6[5327];
@(posedge clk);
#1;data_in = testData6[5328];
@(posedge clk);
#1;data_in = testData6[5329];
@(posedge clk);
#1;data_in = testData6[5330];
@(posedge clk);
#1;data_in = testData6[5331];
@(posedge clk);
#1;data_in = testData6[5332];
@(posedge clk);
#1;data_in = testData6[5333];
@(posedge clk);
#1;data_in = testData6[5334];
@(posedge clk);
#1;data_in = testData6[5335];
@(posedge clk);
#1;data_in = testData6[5336];
@(posedge clk);
#1;data_in = testData6[5337];
@(posedge clk);
#1;data_in = testData6[5338];
@(posedge clk);
#1;data_in = testData6[5339];
@(posedge clk);
#1;data_in = testData6[5340];
@(posedge clk);
#1;data_in = testData6[5341];
@(posedge clk);
#1;data_in = testData6[5342];
@(posedge clk);
#1;data_in = testData6[5343];
@(posedge clk);
#1;data_in = testData6[5344];
@(posedge clk);
#1;data_in = testData6[5345];
@(posedge clk);
#1;data_in = testData6[5346];
@(posedge clk);
#1;data_in = testData6[5347];
@(posedge clk);
#1;data_in = testData6[5348];
@(posedge clk);
#1;data_in = testData6[5349];
@(posedge clk);
#1;data_in = testData6[5350];
@(posedge clk);
#1;data_in = testData6[5351];
@(posedge clk);
#1;data_in = testData6[5352];
@(posedge clk);
#1;data_in = testData6[5353];
@(posedge clk);
#1;data_in = testData6[5354];
@(posedge clk);
#1;data_in = testData6[5355];
@(posedge clk);
#1;data_in = testData6[5356];
@(posedge clk);
#1;data_in = testData6[5357];
@(posedge clk);
#1;data_in = testData6[5358];
@(posedge clk);
#1;data_in = testData6[5359];
@(posedge clk);
#1;data_in = testData6[5360];
@(posedge clk);
#1;data_in = testData6[5361];
@(posedge clk);
#1;data_in = testData6[5362];
@(posedge clk);
#1;data_in = testData6[5363];
@(posedge clk);
#1;data_in = testData6[5364];
@(posedge clk);
#1;data_in = testData6[5365];
@(posedge clk);
#1;data_in = testData6[5366];
@(posedge clk);
#1;data_in = testData6[5367];
@(posedge clk);
#1;data_in = testData6[5368];
@(posedge clk);
#1;data_in = testData6[5369];
@(posedge clk);
#1;data_in = testData6[5370];
@(posedge clk);
#1;data_in = testData6[5371];
@(posedge clk);
#1;data_in = testData6[5372];
@(posedge clk);
#1;data_in = testData6[5373];
@(posedge clk);
#1;data_in = testData6[5374];
@(posedge clk);
#1;data_in = testData6[5375];
@(posedge clk);
#1;data_in = testData6[5376];
@(posedge clk);
#1;data_in = testData6[5377];
@(posedge clk);
#1;data_in = testData6[5378];
@(posedge clk);
#1;data_in = testData6[5379];
@(posedge clk);
#1;data_in = testData6[5380];
@(posedge clk);
#1;data_in = testData6[5381];
@(posedge clk);
#1;data_in = testData6[5382];
@(posedge clk);
#1;data_in = testData6[5383];
@(posedge clk);
#1;data_in = testData6[5384];
@(posedge clk);
#1;data_in = testData6[5385];
@(posedge clk);
#1;data_in = testData6[5386];
@(posedge clk);
#1;data_in = testData6[5387];
@(posedge clk);
#1;data_in = testData6[5388];
@(posedge clk);
#1;data_in = testData6[5389];
@(posedge clk);
#1;data_in = testData6[5390];
@(posedge clk);
#1;data_in = testData6[5391];
@(posedge clk);
#1;data_in = testData6[5392];
@(posedge clk);
#1;data_in = testData6[5393];
@(posedge clk);
#1;data_in = testData6[5394];
@(posedge clk);
#1;data_in = testData6[5395];
@(posedge clk);
#1;data_in = testData6[5396];
@(posedge clk);
#1;data_in = testData6[5397];
@(posedge clk);
#1;data_in = testData6[5398];
@(posedge clk);
#1;data_in = testData6[5399];
@(posedge clk);
#1;data_in = testData6[5400];
@(posedge clk);
#1;data_in = testData6[5401];
@(posedge clk);
#1;data_in = testData6[5402];
@(posedge clk);
#1;data_in = testData6[5403];
@(posedge clk);
#1;data_in = testData6[5404];
@(posedge clk);
#1;data_in = testData6[5405];
@(posedge clk);
#1;data_in = testData6[5406];
@(posedge clk);
#1;data_in = testData6[5407];
@(posedge clk);
#1;data_in = testData6[5408];
@(posedge clk);
#1;data_in = testData6[5409];
@(posedge clk);
#1;data_in = testData6[5410];
@(posedge clk);
#1;data_in = testData6[5411];
@(posedge clk);
#1;data_in = testData6[5412];
@(posedge clk);
#1;data_in = testData6[5413];
@(posedge clk);
#1;data_in = testData6[5414];
@(posedge clk);
#1;data_in = testData6[5415];
@(posedge clk);
#1;data_in = testData6[5416];
@(posedge clk);
#1;data_in = testData6[5417];
@(posedge clk);
#1;data_in = testData6[5418];
@(posedge clk);
#1;data_in = testData6[5419];
@(posedge clk);
#1;data_in = testData6[5420];
@(posedge clk);
#1;data_in = testData6[5421];
@(posedge clk);
#1;data_in = testData6[5422];
@(posedge clk);
#1;data_in = testData6[5423];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[5424]; 
@(posedge clk);
#1;data_in = testData6[5425];
@(posedge clk);
#1;data_in = testData6[5426];
@(posedge clk);
#1;data_in = testData6[5427];
@(posedge clk);
#1;data_in = testData6[5428];
@(posedge clk);
#1;data_in = testData6[5429];
@(posedge clk);
#1;data_in = testData6[5430];
@(posedge clk);
#1;data_in = testData6[5431];
@(posedge clk);
#1;data_in = testData6[5432];
@(posedge clk);
#1;data_in = testData6[5433];
@(posedge clk);
#1;data_in = testData6[5434];
@(posedge clk);
#1;data_in = testData6[5435];
@(posedge clk);
#1;data_in = testData6[5436];
@(posedge clk);
#1;data_in = testData6[5437];
@(posedge clk);
#1;data_in = testData6[5438];
@(posedge clk);
#1;data_in = testData6[5439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[5440];
@(posedge clk);
#1;data_in = testData6[5441];
@(posedge clk);
#1;data_in = testData6[5442];
@(posedge clk);
#1;data_in = testData6[5443];
@(posedge clk);
#1;data_in = testData6[5444];
@(posedge clk);
#1;data_in = testData6[5445];
@(posedge clk);
#1;data_in = testData6[5446];
@(posedge clk);
#1;data_in = testData6[5447];
@(posedge clk);
#1;data_in = testData6[5448];
@(posedge clk);
#1;data_in = testData6[5449];
@(posedge clk);
#1;data_in = testData6[5450];
@(posedge clk);
#1;data_in = testData6[5451];
@(posedge clk);
#1;data_in = testData6[5452];
@(posedge clk);
#1;data_in = testData6[5453];
@(posedge clk);
#1;data_in = testData6[5454];
@(posedge clk);
#1;data_in = testData6[5455];
@(posedge clk);
#1;data_in = testData6[5456];
@(posedge clk);
#1;data_in = testData6[5457];
@(posedge clk);
#1;data_in = testData6[5458];
@(posedge clk);
#1;data_in = testData6[5459];
@(posedge clk);
#1;data_in = testData6[5460];
@(posedge clk);
#1;data_in = testData6[5461];
@(posedge clk);
#1;data_in = testData6[5462];
@(posedge clk);
#1;data_in = testData6[5463];
@(posedge clk);
#1;data_in = testData6[5464];
@(posedge clk);
#1;data_in = testData6[5465];
@(posedge clk);
#1;data_in = testData6[5466];
@(posedge clk);
#1;data_in = testData6[5467];
@(posedge clk);
#1;data_in = testData6[5468];
@(posedge clk);
#1;data_in = testData6[5469];
@(posedge clk);
#1;data_in = testData6[5470];
@(posedge clk);
#1;data_in = testData6[5471];
@(posedge clk);
#1;data_in = testData6[5472];
@(posedge clk);
#1;data_in = testData6[5473];
@(posedge clk);
#1;data_in = testData6[5474];
@(posedge clk);
#1;data_in = testData6[5475];
@(posedge clk);
#1;data_in = testData6[5476];
@(posedge clk);
#1;data_in = testData6[5477];
@(posedge clk);
#1;data_in = testData6[5478];
@(posedge clk);
#1;data_in = testData6[5479];
@(posedge clk);
#1;data_in = testData6[5480];
@(posedge clk);
#1;data_in = testData6[5481];
@(posedge clk);
#1;data_in = testData6[5482];
@(posedge clk);
#1;data_in = testData6[5483];
@(posedge clk);
#1;data_in = testData6[5484];
@(posedge clk);
#1;data_in = testData6[5485];
@(posedge clk);
#1;data_in = testData6[5486];
@(posedge clk);
#1;data_in = testData6[5487];
@(posedge clk);
#1;data_in = testData6[5488];
@(posedge clk);
#1;data_in = testData6[5489];
@(posedge clk);
#1;data_in = testData6[5490];
@(posedge clk);
#1;data_in = testData6[5491];
@(posedge clk);
#1;data_in = testData6[5492];
@(posedge clk);
#1;data_in = testData6[5493];
@(posedge clk);
#1;data_in = testData6[5494];
@(posedge clk);
#1;data_in = testData6[5495];
@(posedge clk);
#1;data_in = testData6[5496];
@(posedge clk);
#1;data_in = testData6[5497];
@(posedge clk);
#1;data_in = testData6[5498];
@(posedge clk);
#1;data_in = testData6[5499];
@(posedge clk);
#1;data_in = testData6[5500];
@(posedge clk);
#1;data_in = testData6[5501];
@(posedge clk);
#1;data_in = testData6[5502];
@(posedge clk);
#1;data_in = testData6[5503];
@(posedge clk);
#1;data_in = testData6[5504];
@(posedge clk);
#1;data_in = testData6[5505];
@(posedge clk);
#1;data_in = testData6[5506];
@(posedge clk);
#1;data_in = testData6[5507];
@(posedge clk);
#1;data_in = testData6[5508];
@(posedge clk);
#1;data_in = testData6[5509];
@(posedge clk);
#1;data_in = testData6[5510];
@(posedge clk);
#1;data_in = testData6[5511];
@(posedge clk);
#1;data_in = testData6[5512];
@(posedge clk);
#1;data_in = testData6[5513];
@(posedge clk);
#1;data_in = testData6[5514];
@(posedge clk);
#1;data_in = testData6[5515];
@(posedge clk);
#1;data_in = testData6[5516];
@(posedge clk);
#1;data_in = testData6[5517];
@(posedge clk);
#1;data_in = testData6[5518];
@(posedge clk);
#1;data_in = testData6[5519];
@(posedge clk);
#1;data_in = testData6[5520];
@(posedge clk);
#1;data_in = testData6[5521];
@(posedge clk);
#1;data_in = testData6[5522];
@(posedge clk);
#1;data_in = testData6[5523];
@(posedge clk);
#1;data_in = testData6[5524];
@(posedge clk);
#1;data_in = testData6[5525];
@(posedge clk);
#1;data_in = testData6[5526];
@(posedge clk);
#1;data_in = testData6[5527];
@(posedge clk);
#1;data_in = testData6[5528];
@(posedge clk);
#1;data_in = testData6[5529];
@(posedge clk);
#1;data_in = testData6[5530];
@(posedge clk);
#1;data_in = testData6[5531];
@(posedge clk);
#1;data_in = testData6[5532];
@(posedge clk);
#1;data_in = testData6[5533];
@(posedge clk);
#1;data_in = testData6[5534];
@(posedge clk);
#1;data_in = testData6[5535];
@(posedge clk);
#1;data_in = testData6[5536];
@(posedge clk);
#1;data_in = testData6[5537];
@(posedge clk);
#1;data_in = testData6[5538];
@(posedge clk);
#1;data_in = testData6[5539];
@(posedge clk);
#1;data_in = testData6[5540];
@(posedge clk);
#1;data_in = testData6[5541];
@(posedge clk);
#1;data_in = testData6[5542];
@(posedge clk);
#1;data_in = testData6[5543];
@(posedge clk);
#1;data_in = testData6[5544];
@(posedge clk);
#1;data_in = testData6[5545];
@(posedge clk);
#1;data_in = testData6[5546];
@(posedge clk);
#1;data_in = testData6[5547];
@(posedge clk);
#1;data_in = testData6[5548];
@(posedge clk);
#1;data_in = testData6[5549];
@(posedge clk);
#1;data_in = testData6[5550];
@(posedge clk);
#1;data_in = testData6[5551];
@(posedge clk);
#1;data_in = testData6[5552];
@(posedge clk);
#1;data_in = testData6[5553];
@(posedge clk);
#1;data_in = testData6[5554];
@(posedge clk);
#1;data_in = testData6[5555];
@(posedge clk);
#1;data_in = testData6[5556];
@(posedge clk);
#1;data_in = testData6[5557];
@(posedge clk);
#1;data_in = testData6[5558];
@(posedge clk);
#1;data_in = testData6[5559];
@(posedge clk);
#1;data_in = testData6[5560];
@(posedge clk);
#1;data_in = testData6[5561];
@(posedge clk);
#1;data_in = testData6[5562];
@(posedge clk);
#1;data_in = testData6[5563];
@(posedge clk);
#1;data_in = testData6[5564];
@(posedge clk);
#1;data_in = testData6[5565];
@(posedge clk);
#1;data_in = testData6[5566];
@(posedge clk);
#1;data_in = testData6[5567];
@(posedge clk);
#1;data_in = testData6[5568];
@(posedge clk);
#1;data_in = testData6[5569];
@(posedge clk);
#1;data_in = testData6[5570];
@(posedge clk);
#1;data_in = testData6[5571];
@(posedge clk);
#1;data_in = testData6[5572];
@(posedge clk);
#1;data_in = testData6[5573];
@(posedge clk);
#1;data_in = testData6[5574];
@(posedge clk);
#1;data_in = testData6[5575];
@(posedge clk);
#1;data_in = testData6[5576];
@(posedge clk);
#1;data_in = testData6[5577];
@(posedge clk);
#1;data_in = testData6[5578];
@(posedge clk);
#1;data_in = testData6[5579];
@(posedge clk);
#1;data_in = testData6[5580];
@(posedge clk);
#1;data_in = testData6[5581];
@(posedge clk);
#1;data_in = testData6[5582];
@(posedge clk);
#1;data_in = testData6[5583];
@(posedge clk);
#1;data_in = testData6[5584];
@(posedge clk);
#1;data_in = testData6[5585];
@(posedge clk);
#1;data_in = testData6[5586];
@(posedge clk);
#1;data_in = testData6[5587];
@(posedge clk);
#1;data_in = testData6[5588];
@(posedge clk);
#1;data_in = testData6[5589];
@(posedge clk);
#1;data_in = testData6[5590];
@(posedge clk);
#1;data_in = testData6[5591];
@(posedge clk);
#1;data_in = testData6[5592];
@(posedge clk);
#1;data_in = testData6[5593];
@(posedge clk);
#1;data_in = testData6[5594];
@(posedge clk);
#1;data_in = testData6[5595];
@(posedge clk);
#1;data_in = testData6[5596];
@(posedge clk);
#1;data_in = testData6[5597];
@(posedge clk);
#1;data_in = testData6[5598];
@(posedge clk);
#1;data_in = testData6[5599];
@(posedge clk);
#1;data_in = testData6[5600];
@(posedge clk);
#1;data_in = testData6[5601];
@(posedge clk);
#1;data_in = testData6[5602];
@(posedge clk);
#1;data_in = testData6[5603];
@(posedge clk);
#1;data_in = testData6[5604];
@(posedge clk);
#1;data_in = testData6[5605];
@(posedge clk);
#1;data_in = testData6[5606];
@(posedge clk);
#1;data_in = testData6[5607];
@(posedge clk);
#1;data_in = testData6[5608];
@(posedge clk);
#1;data_in = testData6[5609];
@(posedge clk);
#1;data_in = testData6[5610];
@(posedge clk);
#1;data_in = testData6[5611];
@(posedge clk);
#1;data_in = testData6[5612];
@(posedge clk);
#1;data_in = testData6[5613];
@(posedge clk);
#1;data_in = testData6[5614];
@(posedge clk);
#1;data_in = testData6[5615];
@(posedge clk);
#1;data_in = testData6[5616];
@(posedge clk);
#1;data_in = testData6[5617];
@(posedge clk);
#1;data_in = testData6[5618];
@(posedge clk);
#1;data_in = testData6[5619];
@(posedge clk);
#1;data_in = testData6[5620];
@(posedge clk);
#1;data_in = testData6[5621];
@(posedge clk);
#1;data_in = testData6[5622];
@(posedge clk);
#1;data_in = testData6[5623];
@(posedge clk);
#1;data_in = testData6[5624];
@(posedge clk);
#1;data_in = testData6[5625];
@(posedge clk);
#1;data_in = testData6[5626];
@(posedge clk);
#1;data_in = testData6[5627];
@(posedge clk);
#1;data_in = testData6[5628];
@(posedge clk);
#1;data_in = testData6[5629];
@(posedge clk);
#1;data_in = testData6[5630];
@(posedge clk);
#1;data_in = testData6[5631];
@(posedge clk);
#1;data_in = testData6[5632];
@(posedge clk);
#1;data_in = testData6[5633];
@(posedge clk);
#1;data_in = testData6[5634];
@(posedge clk);
#1;data_in = testData6[5635];
@(posedge clk);
#1;data_in = testData6[5636];
@(posedge clk);
#1;data_in = testData6[5637];
@(posedge clk);
#1;data_in = testData6[5638];
@(posedge clk);
#1;data_in = testData6[5639];
@(posedge clk);
#1;data_in = testData6[5640];
@(posedge clk);
#1;data_in = testData6[5641];
@(posedge clk);
#1;data_in = testData6[5642];
@(posedge clk);
#1;data_in = testData6[5643];
@(posedge clk);
#1;data_in = testData6[5644];
@(posedge clk);
#1;data_in = testData6[5645];
@(posedge clk);
#1;data_in = testData6[5646];
@(posedge clk);
#1;data_in = testData6[5647];
@(posedge clk);
#1;data_in = testData6[5648];
@(posedge clk);
#1;data_in = testData6[5649];
@(posedge clk);
#1;data_in = testData6[5650];
@(posedge clk);
#1;data_in = testData6[5651];
@(posedge clk);
#1;data_in = testData6[5652];
@(posedge clk);
#1;data_in = testData6[5653];
@(posedge clk);
#1;data_in = testData6[5654];
@(posedge clk);
#1;data_in = testData6[5655];
@(posedge clk);
#1;data_in = testData6[5656];
@(posedge clk);
#1;data_in = testData6[5657];
@(posedge clk);
#1;data_in = testData6[5658];
@(posedge clk);
#1;data_in = testData6[5659];
@(posedge clk);
#1;data_in = testData6[5660];
@(posedge clk);
#1;data_in = testData6[5661];
@(posedge clk);
#1;data_in = testData6[5662];
@(posedge clk);
#1;data_in = testData6[5663];
@(posedge clk);
#1;data_in = testData6[5664];
@(posedge clk);
#1;data_in = testData6[5665];
@(posedge clk);
#1;data_in = testData6[5666];
@(posedge clk);
#1;data_in = testData6[5667];
@(posedge clk);
#1;data_in = testData6[5668];
@(posedge clk);
#1;data_in = testData6[5669];
@(posedge clk);
#1;data_in = testData6[5670];
@(posedge clk);
#1;data_in = testData6[5671];
@(posedge clk);
#1;data_in = testData6[5672];
@(posedge clk);
#1;data_in = testData6[5673];
@(posedge clk);
#1;data_in = testData6[5674];
@(posedge clk);
#1;data_in = testData6[5675];
@(posedge clk);
#1;data_in = testData6[5676];
@(posedge clk);
#1;data_in = testData6[5677];
@(posedge clk);
#1;data_in = testData6[5678];
@(posedge clk);
#1;data_in = testData6[5679];
@(posedge clk);
#1;data_in = testData6[5680];
@(posedge clk);
#1;data_in = testData6[5681];
@(posedge clk);
#1;data_in = testData6[5682];
@(posedge clk);
#1;data_in = testData6[5683];
@(posedge clk);
#1;data_in = testData6[5684];
@(posedge clk);
#1;data_in = testData6[5685];
@(posedge clk);
#1;data_in = testData6[5686];
@(posedge clk);
#1;data_in = testData6[5687];
@(posedge clk);
#1;data_in = testData6[5688];
@(posedge clk);
#1;data_in = testData6[5689];
@(posedge clk);
#1;data_in = testData6[5690];
@(posedge clk);
#1;data_in = testData6[5691];
@(posedge clk);
#1;data_in = testData6[5692];
@(posedge clk);
#1;data_in = testData6[5693];
@(posedge clk);
#1;data_in = testData6[5694];
@(posedge clk);
#1;data_in = testData6[5695];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[5696]; 
@(posedge clk);
#1;data_in = testData6[5697];
@(posedge clk);
#1;data_in = testData6[5698];
@(posedge clk);
#1;data_in = testData6[5699];
@(posedge clk);
#1;data_in = testData6[5700];
@(posedge clk);
#1;data_in = testData6[5701];
@(posedge clk);
#1;data_in = testData6[5702];
@(posedge clk);
#1;data_in = testData6[5703];
@(posedge clk);
#1;data_in = testData6[5704];
@(posedge clk);
#1;data_in = testData6[5705];
@(posedge clk);
#1;data_in = testData6[5706];
@(posedge clk);
#1;data_in = testData6[5707];
@(posedge clk);
#1;data_in = testData6[5708];
@(posedge clk);
#1;data_in = testData6[5709];
@(posedge clk);
#1;data_in = testData6[5710];
@(posedge clk);
#1;data_in = testData6[5711];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[5712];
@(posedge clk);
#1;data_in = testData6[5713];
@(posedge clk);
#1;data_in = testData6[5714];
@(posedge clk);
#1;data_in = testData6[5715];
@(posedge clk);
#1;data_in = testData6[5716];
@(posedge clk);
#1;data_in = testData6[5717];
@(posedge clk);
#1;data_in = testData6[5718];
@(posedge clk);
#1;data_in = testData6[5719];
@(posedge clk);
#1;data_in = testData6[5720];
@(posedge clk);
#1;data_in = testData6[5721];
@(posedge clk);
#1;data_in = testData6[5722];
@(posedge clk);
#1;data_in = testData6[5723];
@(posedge clk);
#1;data_in = testData6[5724];
@(posedge clk);
#1;data_in = testData6[5725];
@(posedge clk);
#1;data_in = testData6[5726];
@(posedge clk);
#1;data_in = testData6[5727];
@(posedge clk);
#1;data_in = testData6[5728];
@(posedge clk);
#1;data_in = testData6[5729];
@(posedge clk);
#1;data_in = testData6[5730];
@(posedge clk);
#1;data_in = testData6[5731];
@(posedge clk);
#1;data_in = testData6[5732];
@(posedge clk);
#1;data_in = testData6[5733];
@(posedge clk);
#1;data_in = testData6[5734];
@(posedge clk);
#1;data_in = testData6[5735];
@(posedge clk);
#1;data_in = testData6[5736];
@(posedge clk);
#1;data_in = testData6[5737];
@(posedge clk);
#1;data_in = testData6[5738];
@(posedge clk);
#1;data_in = testData6[5739];
@(posedge clk);
#1;data_in = testData6[5740];
@(posedge clk);
#1;data_in = testData6[5741];
@(posedge clk);
#1;data_in = testData6[5742];
@(posedge clk);
#1;data_in = testData6[5743];
@(posedge clk);
#1;data_in = testData6[5744];
@(posedge clk);
#1;data_in = testData6[5745];
@(posedge clk);
#1;data_in = testData6[5746];
@(posedge clk);
#1;data_in = testData6[5747];
@(posedge clk);
#1;data_in = testData6[5748];
@(posedge clk);
#1;data_in = testData6[5749];
@(posedge clk);
#1;data_in = testData6[5750];
@(posedge clk);
#1;data_in = testData6[5751];
@(posedge clk);
#1;data_in = testData6[5752];
@(posedge clk);
#1;data_in = testData6[5753];
@(posedge clk);
#1;data_in = testData6[5754];
@(posedge clk);
#1;data_in = testData6[5755];
@(posedge clk);
#1;data_in = testData6[5756];
@(posedge clk);
#1;data_in = testData6[5757];
@(posedge clk);
#1;data_in = testData6[5758];
@(posedge clk);
#1;data_in = testData6[5759];
@(posedge clk);
#1;data_in = testData6[5760];
@(posedge clk);
#1;data_in = testData6[5761];
@(posedge clk);
#1;data_in = testData6[5762];
@(posedge clk);
#1;data_in = testData6[5763];
@(posedge clk);
#1;data_in = testData6[5764];
@(posedge clk);
#1;data_in = testData6[5765];
@(posedge clk);
#1;data_in = testData6[5766];
@(posedge clk);
#1;data_in = testData6[5767];
@(posedge clk);
#1;data_in = testData6[5768];
@(posedge clk);
#1;data_in = testData6[5769];
@(posedge clk);
#1;data_in = testData6[5770];
@(posedge clk);
#1;data_in = testData6[5771];
@(posedge clk);
#1;data_in = testData6[5772];
@(posedge clk);
#1;data_in = testData6[5773];
@(posedge clk);
#1;data_in = testData6[5774];
@(posedge clk);
#1;data_in = testData6[5775];
@(posedge clk);
#1;data_in = testData6[5776];
@(posedge clk);
#1;data_in = testData6[5777];
@(posedge clk);
#1;data_in = testData6[5778];
@(posedge clk);
#1;data_in = testData6[5779];
@(posedge clk);
#1;data_in = testData6[5780];
@(posedge clk);
#1;data_in = testData6[5781];
@(posedge clk);
#1;data_in = testData6[5782];
@(posedge clk);
#1;data_in = testData6[5783];
@(posedge clk);
#1;data_in = testData6[5784];
@(posedge clk);
#1;data_in = testData6[5785];
@(posedge clk);
#1;data_in = testData6[5786];
@(posedge clk);
#1;data_in = testData6[5787];
@(posedge clk);
#1;data_in = testData6[5788];
@(posedge clk);
#1;data_in = testData6[5789];
@(posedge clk);
#1;data_in = testData6[5790];
@(posedge clk);
#1;data_in = testData6[5791];
@(posedge clk);
#1;data_in = testData6[5792];
@(posedge clk);
#1;data_in = testData6[5793];
@(posedge clk);
#1;data_in = testData6[5794];
@(posedge clk);
#1;data_in = testData6[5795];
@(posedge clk);
#1;data_in = testData6[5796];
@(posedge clk);
#1;data_in = testData6[5797];
@(posedge clk);
#1;data_in = testData6[5798];
@(posedge clk);
#1;data_in = testData6[5799];
@(posedge clk);
#1;data_in = testData6[5800];
@(posedge clk);
#1;data_in = testData6[5801];
@(posedge clk);
#1;data_in = testData6[5802];
@(posedge clk);
#1;data_in = testData6[5803];
@(posedge clk);
#1;data_in = testData6[5804];
@(posedge clk);
#1;data_in = testData6[5805];
@(posedge clk);
#1;data_in = testData6[5806];
@(posedge clk);
#1;data_in = testData6[5807];
@(posedge clk);
#1;data_in = testData6[5808];
@(posedge clk);
#1;data_in = testData6[5809];
@(posedge clk);
#1;data_in = testData6[5810];
@(posedge clk);
#1;data_in = testData6[5811];
@(posedge clk);
#1;data_in = testData6[5812];
@(posedge clk);
#1;data_in = testData6[5813];
@(posedge clk);
#1;data_in = testData6[5814];
@(posedge clk);
#1;data_in = testData6[5815];
@(posedge clk);
#1;data_in = testData6[5816];
@(posedge clk);
#1;data_in = testData6[5817];
@(posedge clk);
#1;data_in = testData6[5818];
@(posedge clk);
#1;data_in = testData6[5819];
@(posedge clk);
#1;data_in = testData6[5820];
@(posedge clk);
#1;data_in = testData6[5821];
@(posedge clk);
#1;data_in = testData6[5822];
@(posedge clk);
#1;data_in = testData6[5823];
@(posedge clk);
#1;data_in = testData6[5824];
@(posedge clk);
#1;data_in = testData6[5825];
@(posedge clk);
#1;data_in = testData6[5826];
@(posedge clk);
#1;data_in = testData6[5827];
@(posedge clk);
#1;data_in = testData6[5828];
@(posedge clk);
#1;data_in = testData6[5829];
@(posedge clk);
#1;data_in = testData6[5830];
@(posedge clk);
#1;data_in = testData6[5831];
@(posedge clk);
#1;data_in = testData6[5832];
@(posedge clk);
#1;data_in = testData6[5833];
@(posedge clk);
#1;data_in = testData6[5834];
@(posedge clk);
#1;data_in = testData6[5835];
@(posedge clk);
#1;data_in = testData6[5836];
@(posedge clk);
#1;data_in = testData6[5837];
@(posedge clk);
#1;data_in = testData6[5838];
@(posedge clk);
#1;data_in = testData6[5839];
@(posedge clk);
#1;data_in = testData6[5840];
@(posedge clk);
#1;data_in = testData6[5841];
@(posedge clk);
#1;data_in = testData6[5842];
@(posedge clk);
#1;data_in = testData6[5843];
@(posedge clk);
#1;data_in = testData6[5844];
@(posedge clk);
#1;data_in = testData6[5845];
@(posedge clk);
#1;data_in = testData6[5846];
@(posedge clk);
#1;data_in = testData6[5847];
@(posedge clk);
#1;data_in = testData6[5848];
@(posedge clk);
#1;data_in = testData6[5849];
@(posedge clk);
#1;data_in = testData6[5850];
@(posedge clk);
#1;data_in = testData6[5851];
@(posedge clk);
#1;data_in = testData6[5852];
@(posedge clk);
#1;data_in = testData6[5853];
@(posedge clk);
#1;data_in = testData6[5854];
@(posedge clk);
#1;data_in = testData6[5855];
@(posedge clk);
#1;data_in = testData6[5856];
@(posedge clk);
#1;data_in = testData6[5857];
@(posedge clk);
#1;data_in = testData6[5858];
@(posedge clk);
#1;data_in = testData6[5859];
@(posedge clk);
#1;data_in = testData6[5860];
@(posedge clk);
#1;data_in = testData6[5861];
@(posedge clk);
#1;data_in = testData6[5862];
@(posedge clk);
#1;data_in = testData6[5863];
@(posedge clk);
#1;data_in = testData6[5864];
@(posedge clk);
#1;data_in = testData6[5865];
@(posedge clk);
#1;data_in = testData6[5866];
@(posedge clk);
#1;data_in = testData6[5867];
@(posedge clk);
#1;data_in = testData6[5868];
@(posedge clk);
#1;data_in = testData6[5869];
@(posedge clk);
#1;data_in = testData6[5870];
@(posedge clk);
#1;data_in = testData6[5871];
@(posedge clk);
#1;data_in = testData6[5872];
@(posedge clk);
#1;data_in = testData6[5873];
@(posedge clk);
#1;data_in = testData6[5874];
@(posedge clk);
#1;data_in = testData6[5875];
@(posedge clk);
#1;data_in = testData6[5876];
@(posedge clk);
#1;data_in = testData6[5877];
@(posedge clk);
#1;data_in = testData6[5878];
@(posedge clk);
#1;data_in = testData6[5879];
@(posedge clk);
#1;data_in = testData6[5880];
@(posedge clk);
#1;data_in = testData6[5881];
@(posedge clk);
#1;data_in = testData6[5882];
@(posedge clk);
#1;data_in = testData6[5883];
@(posedge clk);
#1;data_in = testData6[5884];
@(posedge clk);
#1;data_in = testData6[5885];
@(posedge clk);
#1;data_in = testData6[5886];
@(posedge clk);
#1;data_in = testData6[5887];
@(posedge clk);
#1;data_in = testData6[5888];
@(posedge clk);
#1;data_in = testData6[5889];
@(posedge clk);
#1;data_in = testData6[5890];
@(posedge clk);
#1;data_in = testData6[5891];
@(posedge clk);
#1;data_in = testData6[5892];
@(posedge clk);
#1;data_in = testData6[5893];
@(posedge clk);
#1;data_in = testData6[5894];
@(posedge clk);
#1;data_in = testData6[5895];
@(posedge clk);
#1;data_in = testData6[5896];
@(posedge clk);
#1;data_in = testData6[5897];
@(posedge clk);
#1;data_in = testData6[5898];
@(posedge clk);
#1;data_in = testData6[5899];
@(posedge clk);
#1;data_in = testData6[5900];
@(posedge clk);
#1;data_in = testData6[5901];
@(posedge clk);
#1;data_in = testData6[5902];
@(posedge clk);
#1;data_in = testData6[5903];
@(posedge clk);
#1;data_in = testData6[5904];
@(posedge clk);
#1;data_in = testData6[5905];
@(posedge clk);
#1;data_in = testData6[5906];
@(posedge clk);
#1;data_in = testData6[5907];
@(posedge clk);
#1;data_in = testData6[5908];
@(posedge clk);
#1;data_in = testData6[5909];
@(posedge clk);
#1;data_in = testData6[5910];
@(posedge clk);
#1;data_in = testData6[5911];
@(posedge clk);
#1;data_in = testData6[5912];
@(posedge clk);
#1;data_in = testData6[5913];
@(posedge clk);
#1;data_in = testData6[5914];
@(posedge clk);
#1;data_in = testData6[5915];
@(posedge clk);
#1;data_in = testData6[5916];
@(posedge clk);
#1;data_in = testData6[5917];
@(posedge clk);
#1;data_in = testData6[5918];
@(posedge clk);
#1;data_in = testData6[5919];
@(posedge clk);
#1;data_in = testData6[5920];
@(posedge clk);
#1;data_in = testData6[5921];
@(posedge clk);
#1;data_in = testData6[5922];
@(posedge clk);
#1;data_in = testData6[5923];
@(posedge clk);
#1;data_in = testData6[5924];
@(posedge clk);
#1;data_in = testData6[5925];
@(posedge clk);
#1;data_in = testData6[5926];
@(posedge clk);
#1;data_in = testData6[5927];
@(posedge clk);
#1;data_in = testData6[5928];
@(posedge clk);
#1;data_in = testData6[5929];
@(posedge clk);
#1;data_in = testData6[5930];
@(posedge clk);
#1;data_in = testData6[5931];
@(posedge clk);
#1;data_in = testData6[5932];
@(posedge clk);
#1;data_in = testData6[5933];
@(posedge clk);
#1;data_in = testData6[5934];
@(posedge clk);
#1;data_in = testData6[5935];
@(posedge clk);
#1;data_in = testData6[5936];
@(posedge clk);
#1;data_in = testData6[5937];
@(posedge clk);
#1;data_in = testData6[5938];
@(posedge clk);
#1;data_in = testData6[5939];
@(posedge clk);
#1;data_in = testData6[5940];
@(posedge clk);
#1;data_in = testData6[5941];
@(posedge clk);
#1;data_in = testData6[5942];
@(posedge clk);
#1;data_in = testData6[5943];
@(posedge clk);
#1;data_in = testData6[5944];
@(posedge clk);
#1;data_in = testData6[5945];
@(posedge clk);
#1;data_in = testData6[5946];
@(posedge clk);
#1;data_in = testData6[5947];
@(posedge clk);
#1;data_in = testData6[5948];
@(posedge clk);
#1;data_in = testData6[5949];
@(posedge clk);
#1;data_in = testData6[5950];
@(posedge clk);
#1;data_in = testData6[5951];
@(posedge clk);
#1;data_in = testData6[5952];
@(posedge clk);
#1;data_in = testData6[5953];
@(posedge clk);
#1;data_in = testData6[5954];
@(posedge clk);
#1;data_in = testData6[5955];
@(posedge clk);
#1;data_in = testData6[5956];
@(posedge clk);
#1;data_in = testData6[5957];
@(posedge clk);
#1;data_in = testData6[5958];
@(posedge clk);
#1;data_in = testData6[5959];
@(posedge clk);
#1;data_in = testData6[5960];
@(posedge clk);
#1;data_in = testData6[5961];
@(posedge clk);
#1;data_in = testData6[5962];
@(posedge clk);
#1;data_in = testData6[5963];
@(posedge clk);
#1;data_in = testData6[5964];
@(posedge clk);
#1;data_in = testData6[5965];
@(posedge clk);
#1;data_in = testData6[5966];
@(posedge clk);
#1;data_in = testData6[5967];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[5968]; 
@(posedge clk);
#1;data_in = testData6[5969];
@(posedge clk);
#1;data_in = testData6[5970];
@(posedge clk);
#1;data_in = testData6[5971];
@(posedge clk);
#1;data_in = testData6[5972];
@(posedge clk);
#1;data_in = testData6[5973];
@(posedge clk);
#1;data_in = testData6[5974];
@(posedge clk);
#1;data_in = testData6[5975];
@(posedge clk);
#1;data_in = testData6[5976];
@(posedge clk);
#1;data_in = testData6[5977];
@(posedge clk);
#1;data_in = testData6[5978];
@(posedge clk);
#1;data_in = testData6[5979];
@(posedge clk);
#1;data_in = testData6[5980];
@(posedge clk);
#1;data_in = testData6[5981];
@(posedge clk);
#1;data_in = testData6[5982];
@(posedge clk);
#1;data_in = testData6[5983];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[5984];
@(posedge clk);
#1;data_in = testData6[5985];
@(posedge clk);
#1;data_in = testData6[5986];
@(posedge clk);
#1;data_in = testData6[5987];
@(posedge clk);
#1;data_in = testData6[5988];
@(posedge clk);
#1;data_in = testData6[5989];
@(posedge clk);
#1;data_in = testData6[5990];
@(posedge clk);
#1;data_in = testData6[5991];
@(posedge clk);
#1;data_in = testData6[5992];
@(posedge clk);
#1;data_in = testData6[5993];
@(posedge clk);
#1;data_in = testData6[5994];
@(posedge clk);
#1;data_in = testData6[5995];
@(posedge clk);
#1;data_in = testData6[5996];
@(posedge clk);
#1;data_in = testData6[5997];
@(posedge clk);
#1;data_in = testData6[5998];
@(posedge clk);
#1;data_in = testData6[5999];
@(posedge clk);
#1;data_in = testData6[6000];
@(posedge clk);
#1;data_in = testData6[6001];
@(posedge clk);
#1;data_in = testData6[6002];
@(posedge clk);
#1;data_in = testData6[6003];
@(posedge clk);
#1;data_in = testData6[6004];
@(posedge clk);
#1;data_in = testData6[6005];
@(posedge clk);
#1;data_in = testData6[6006];
@(posedge clk);
#1;data_in = testData6[6007];
@(posedge clk);
#1;data_in = testData6[6008];
@(posedge clk);
#1;data_in = testData6[6009];
@(posedge clk);
#1;data_in = testData6[6010];
@(posedge clk);
#1;data_in = testData6[6011];
@(posedge clk);
#1;data_in = testData6[6012];
@(posedge clk);
#1;data_in = testData6[6013];
@(posedge clk);
#1;data_in = testData6[6014];
@(posedge clk);
#1;data_in = testData6[6015];
@(posedge clk);
#1;data_in = testData6[6016];
@(posedge clk);
#1;data_in = testData6[6017];
@(posedge clk);
#1;data_in = testData6[6018];
@(posedge clk);
#1;data_in = testData6[6019];
@(posedge clk);
#1;data_in = testData6[6020];
@(posedge clk);
#1;data_in = testData6[6021];
@(posedge clk);
#1;data_in = testData6[6022];
@(posedge clk);
#1;data_in = testData6[6023];
@(posedge clk);
#1;data_in = testData6[6024];
@(posedge clk);
#1;data_in = testData6[6025];
@(posedge clk);
#1;data_in = testData6[6026];
@(posedge clk);
#1;data_in = testData6[6027];
@(posedge clk);
#1;data_in = testData6[6028];
@(posedge clk);
#1;data_in = testData6[6029];
@(posedge clk);
#1;data_in = testData6[6030];
@(posedge clk);
#1;data_in = testData6[6031];
@(posedge clk);
#1;data_in = testData6[6032];
@(posedge clk);
#1;data_in = testData6[6033];
@(posedge clk);
#1;data_in = testData6[6034];
@(posedge clk);
#1;data_in = testData6[6035];
@(posedge clk);
#1;data_in = testData6[6036];
@(posedge clk);
#1;data_in = testData6[6037];
@(posedge clk);
#1;data_in = testData6[6038];
@(posedge clk);
#1;data_in = testData6[6039];
@(posedge clk);
#1;data_in = testData6[6040];
@(posedge clk);
#1;data_in = testData6[6041];
@(posedge clk);
#1;data_in = testData6[6042];
@(posedge clk);
#1;data_in = testData6[6043];
@(posedge clk);
#1;data_in = testData6[6044];
@(posedge clk);
#1;data_in = testData6[6045];
@(posedge clk);
#1;data_in = testData6[6046];
@(posedge clk);
#1;data_in = testData6[6047];
@(posedge clk);
#1;data_in = testData6[6048];
@(posedge clk);
#1;data_in = testData6[6049];
@(posedge clk);
#1;data_in = testData6[6050];
@(posedge clk);
#1;data_in = testData6[6051];
@(posedge clk);
#1;data_in = testData6[6052];
@(posedge clk);
#1;data_in = testData6[6053];
@(posedge clk);
#1;data_in = testData6[6054];
@(posedge clk);
#1;data_in = testData6[6055];
@(posedge clk);
#1;data_in = testData6[6056];
@(posedge clk);
#1;data_in = testData6[6057];
@(posedge clk);
#1;data_in = testData6[6058];
@(posedge clk);
#1;data_in = testData6[6059];
@(posedge clk);
#1;data_in = testData6[6060];
@(posedge clk);
#1;data_in = testData6[6061];
@(posedge clk);
#1;data_in = testData6[6062];
@(posedge clk);
#1;data_in = testData6[6063];
@(posedge clk);
#1;data_in = testData6[6064];
@(posedge clk);
#1;data_in = testData6[6065];
@(posedge clk);
#1;data_in = testData6[6066];
@(posedge clk);
#1;data_in = testData6[6067];
@(posedge clk);
#1;data_in = testData6[6068];
@(posedge clk);
#1;data_in = testData6[6069];
@(posedge clk);
#1;data_in = testData6[6070];
@(posedge clk);
#1;data_in = testData6[6071];
@(posedge clk);
#1;data_in = testData6[6072];
@(posedge clk);
#1;data_in = testData6[6073];
@(posedge clk);
#1;data_in = testData6[6074];
@(posedge clk);
#1;data_in = testData6[6075];
@(posedge clk);
#1;data_in = testData6[6076];
@(posedge clk);
#1;data_in = testData6[6077];
@(posedge clk);
#1;data_in = testData6[6078];
@(posedge clk);
#1;data_in = testData6[6079];
@(posedge clk);
#1;data_in = testData6[6080];
@(posedge clk);
#1;data_in = testData6[6081];
@(posedge clk);
#1;data_in = testData6[6082];
@(posedge clk);
#1;data_in = testData6[6083];
@(posedge clk);
#1;data_in = testData6[6084];
@(posedge clk);
#1;data_in = testData6[6085];
@(posedge clk);
#1;data_in = testData6[6086];
@(posedge clk);
#1;data_in = testData6[6087];
@(posedge clk);
#1;data_in = testData6[6088];
@(posedge clk);
#1;data_in = testData6[6089];
@(posedge clk);
#1;data_in = testData6[6090];
@(posedge clk);
#1;data_in = testData6[6091];
@(posedge clk);
#1;data_in = testData6[6092];
@(posedge clk);
#1;data_in = testData6[6093];
@(posedge clk);
#1;data_in = testData6[6094];
@(posedge clk);
#1;data_in = testData6[6095];
@(posedge clk);
#1;data_in = testData6[6096];
@(posedge clk);
#1;data_in = testData6[6097];
@(posedge clk);
#1;data_in = testData6[6098];
@(posedge clk);
#1;data_in = testData6[6099];
@(posedge clk);
#1;data_in = testData6[6100];
@(posedge clk);
#1;data_in = testData6[6101];
@(posedge clk);
#1;data_in = testData6[6102];
@(posedge clk);
#1;data_in = testData6[6103];
@(posedge clk);
#1;data_in = testData6[6104];
@(posedge clk);
#1;data_in = testData6[6105];
@(posedge clk);
#1;data_in = testData6[6106];
@(posedge clk);
#1;data_in = testData6[6107];
@(posedge clk);
#1;data_in = testData6[6108];
@(posedge clk);
#1;data_in = testData6[6109];
@(posedge clk);
#1;data_in = testData6[6110];
@(posedge clk);
#1;data_in = testData6[6111];
@(posedge clk);
#1;data_in = testData6[6112];
@(posedge clk);
#1;data_in = testData6[6113];
@(posedge clk);
#1;data_in = testData6[6114];
@(posedge clk);
#1;data_in = testData6[6115];
@(posedge clk);
#1;data_in = testData6[6116];
@(posedge clk);
#1;data_in = testData6[6117];
@(posedge clk);
#1;data_in = testData6[6118];
@(posedge clk);
#1;data_in = testData6[6119];
@(posedge clk);
#1;data_in = testData6[6120];
@(posedge clk);
#1;data_in = testData6[6121];
@(posedge clk);
#1;data_in = testData6[6122];
@(posedge clk);
#1;data_in = testData6[6123];
@(posedge clk);
#1;data_in = testData6[6124];
@(posedge clk);
#1;data_in = testData6[6125];
@(posedge clk);
#1;data_in = testData6[6126];
@(posedge clk);
#1;data_in = testData6[6127];
@(posedge clk);
#1;data_in = testData6[6128];
@(posedge clk);
#1;data_in = testData6[6129];
@(posedge clk);
#1;data_in = testData6[6130];
@(posedge clk);
#1;data_in = testData6[6131];
@(posedge clk);
#1;data_in = testData6[6132];
@(posedge clk);
#1;data_in = testData6[6133];
@(posedge clk);
#1;data_in = testData6[6134];
@(posedge clk);
#1;data_in = testData6[6135];
@(posedge clk);
#1;data_in = testData6[6136];
@(posedge clk);
#1;data_in = testData6[6137];
@(posedge clk);
#1;data_in = testData6[6138];
@(posedge clk);
#1;data_in = testData6[6139];
@(posedge clk);
#1;data_in = testData6[6140];
@(posedge clk);
#1;data_in = testData6[6141];
@(posedge clk);
#1;data_in = testData6[6142];
@(posedge clk);
#1;data_in = testData6[6143];
@(posedge clk);
#1;data_in = testData6[6144];
@(posedge clk);
#1;data_in = testData6[6145];
@(posedge clk);
#1;data_in = testData6[6146];
@(posedge clk);
#1;data_in = testData6[6147];
@(posedge clk);
#1;data_in = testData6[6148];
@(posedge clk);
#1;data_in = testData6[6149];
@(posedge clk);
#1;data_in = testData6[6150];
@(posedge clk);
#1;data_in = testData6[6151];
@(posedge clk);
#1;data_in = testData6[6152];
@(posedge clk);
#1;data_in = testData6[6153];
@(posedge clk);
#1;data_in = testData6[6154];
@(posedge clk);
#1;data_in = testData6[6155];
@(posedge clk);
#1;data_in = testData6[6156];
@(posedge clk);
#1;data_in = testData6[6157];
@(posedge clk);
#1;data_in = testData6[6158];
@(posedge clk);
#1;data_in = testData6[6159];
@(posedge clk);
#1;data_in = testData6[6160];
@(posedge clk);
#1;data_in = testData6[6161];
@(posedge clk);
#1;data_in = testData6[6162];
@(posedge clk);
#1;data_in = testData6[6163];
@(posedge clk);
#1;data_in = testData6[6164];
@(posedge clk);
#1;data_in = testData6[6165];
@(posedge clk);
#1;data_in = testData6[6166];
@(posedge clk);
#1;data_in = testData6[6167];
@(posedge clk);
#1;data_in = testData6[6168];
@(posedge clk);
#1;data_in = testData6[6169];
@(posedge clk);
#1;data_in = testData6[6170];
@(posedge clk);
#1;data_in = testData6[6171];
@(posedge clk);
#1;data_in = testData6[6172];
@(posedge clk);
#1;data_in = testData6[6173];
@(posedge clk);
#1;data_in = testData6[6174];
@(posedge clk);
#1;data_in = testData6[6175];
@(posedge clk);
#1;data_in = testData6[6176];
@(posedge clk);
#1;data_in = testData6[6177];
@(posedge clk);
#1;data_in = testData6[6178];
@(posedge clk);
#1;data_in = testData6[6179];
@(posedge clk);
#1;data_in = testData6[6180];
@(posedge clk);
#1;data_in = testData6[6181];
@(posedge clk);
#1;data_in = testData6[6182];
@(posedge clk);
#1;data_in = testData6[6183];
@(posedge clk);
#1;data_in = testData6[6184];
@(posedge clk);
#1;data_in = testData6[6185];
@(posedge clk);
#1;data_in = testData6[6186];
@(posedge clk);
#1;data_in = testData6[6187];
@(posedge clk);
#1;data_in = testData6[6188];
@(posedge clk);
#1;data_in = testData6[6189];
@(posedge clk);
#1;data_in = testData6[6190];
@(posedge clk);
#1;data_in = testData6[6191];
@(posedge clk);
#1;data_in = testData6[6192];
@(posedge clk);
#1;data_in = testData6[6193];
@(posedge clk);
#1;data_in = testData6[6194];
@(posedge clk);
#1;data_in = testData6[6195];
@(posedge clk);
#1;data_in = testData6[6196];
@(posedge clk);
#1;data_in = testData6[6197];
@(posedge clk);
#1;data_in = testData6[6198];
@(posedge clk);
#1;data_in = testData6[6199];
@(posedge clk);
#1;data_in = testData6[6200];
@(posedge clk);
#1;data_in = testData6[6201];
@(posedge clk);
#1;data_in = testData6[6202];
@(posedge clk);
#1;data_in = testData6[6203];
@(posedge clk);
#1;data_in = testData6[6204];
@(posedge clk);
#1;data_in = testData6[6205];
@(posedge clk);
#1;data_in = testData6[6206];
@(posedge clk);
#1;data_in = testData6[6207];
@(posedge clk);
#1;data_in = testData6[6208];
@(posedge clk);
#1;data_in = testData6[6209];
@(posedge clk);
#1;data_in = testData6[6210];
@(posedge clk);
#1;data_in = testData6[6211];
@(posedge clk);
#1;data_in = testData6[6212];
@(posedge clk);
#1;data_in = testData6[6213];
@(posedge clk);
#1;data_in = testData6[6214];
@(posedge clk);
#1;data_in = testData6[6215];
@(posedge clk);
#1;data_in = testData6[6216];
@(posedge clk);
#1;data_in = testData6[6217];
@(posedge clk);
#1;data_in = testData6[6218];
@(posedge clk);
#1;data_in = testData6[6219];
@(posedge clk);
#1;data_in = testData6[6220];
@(posedge clk);
#1;data_in = testData6[6221];
@(posedge clk);
#1;data_in = testData6[6222];
@(posedge clk);
#1;data_in = testData6[6223];
@(posedge clk);
#1;data_in = testData6[6224];
@(posedge clk);
#1;data_in = testData6[6225];
@(posedge clk);
#1;data_in = testData6[6226];
@(posedge clk);
#1;data_in = testData6[6227];
@(posedge clk);
#1;data_in = testData6[6228];
@(posedge clk);
#1;data_in = testData6[6229];
@(posedge clk);
#1;data_in = testData6[6230];
@(posedge clk);
#1;data_in = testData6[6231];
@(posedge clk);
#1;data_in = testData6[6232];
@(posedge clk);
#1;data_in = testData6[6233];
@(posedge clk);
#1;data_in = testData6[6234];
@(posedge clk);
#1;data_in = testData6[6235];
@(posedge clk);
#1;data_in = testData6[6236];
@(posedge clk);
#1;data_in = testData6[6237];
@(posedge clk);
#1;data_in = testData6[6238];
@(posedge clk);
#1;data_in = testData6[6239];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[6240]; 
@(posedge clk);
#1;data_in = testData6[6241];
@(posedge clk);
#1;data_in = testData6[6242];
@(posedge clk);
#1;data_in = testData6[6243];
@(posedge clk);
#1;data_in = testData6[6244];
@(posedge clk);
#1;data_in = testData6[6245];
@(posedge clk);
#1;data_in = testData6[6246];
@(posedge clk);
#1;data_in = testData6[6247];
@(posedge clk);
#1;data_in = testData6[6248];
@(posedge clk);
#1;data_in = testData6[6249];
@(posedge clk);
#1;data_in = testData6[6250];
@(posedge clk);
#1;data_in = testData6[6251];
@(posedge clk);
#1;data_in = testData6[6252];
@(posedge clk);
#1;data_in = testData6[6253];
@(posedge clk);
#1;data_in = testData6[6254];
@(posedge clk);
#1;data_in = testData6[6255];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[6256];
@(posedge clk);
#1;data_in = testData6[6257];
@(posedge clk);
#1;data_in = testData6[6258];
@(posedge clk);
#1;data_in = testData6[6259];
@(posedge clk);
#1;data_in = testData6[6260];
@(posedge clk);
#1;data_in = testData6[6261];
@(posedge clk);
#1;data_in = testData6[6262];
@(posedge clk);
#1;data_in = testData6[6263];
@(posedge clk);
#1;data_in = testData6[6264];
@(posedge clk);
#1;data_in = testData6[6265];
@(posedge clk);
#1;data_in = testData6[6266];
@(posedge clk);
#1;data_in = testData6[6267];
@(posedge clk);
#1;data_in = testData6[6268];
@(posedge clk);
#1;data_in = testData6[6269];
@(posedge clk);
#1;data_in = testData6[6270];
@(posedge clk);
#1;data_in = testData6[6271];
@(posedge clk);
#1;data_in = testData6[6272];
@(posedge clk);
#1;data_in = testData6[6273];
@(posedge clk);
#1;data_in = testData6[6274];
@(posedge clk);
#1;data_in = testData6[6275];
@(posedge clk);
#1;data_in = testData6[6276];
@(posedge clk);
#1;data_in = testData6[6277];
@(posedge clk);
#1;data_in = testData6[6278];
@(posedge clk);
#1;data_in = testData6[6279];
@(posedge clk);
#1;data_in = testData6[6280];
@(posedge clk);
#1;data_in = testData6[6281];
@(posedge clk);
#1;data_in = testData6[6282];
@(posedge clk);
#1;data_in = testData6[6283];
@(posedge clk);
#1;data_in = testData6[6284];
@(posedge clk);
#1;data_in = testData6[6285];
@(posedge clk);
#1;data_in = testData6[6286];
@(posedge clk);
#1;data_in = testData6[6287];
@(posedge clk);
#1;data_in = testData6[6288];
@(posedge clk);
#1;data_in = testData6[6289];
@(posedge clk);
#1;data_in = testData6[6290];
@(posedge clk);
#1;data_in = testData6[6291];
@(posedge clk);
#1;data_in = testData6[6292];
@(posedge clk);
#1;data_in = testData6[6293];
@(posedge clk);
#1;data_in = testData6[6294];
@(posedge clk);
#1;data_in = testData6[6295];
@(posedge clk);
#1;data_in = testData6[6296];
@(posedge clk);
#1;data_in = testData6[6297];
@(posedge clk);
#1;data_in = testData6[6298];
@(posedge clk);
#1;data_in = testData6[6299];
@(posedge clk);
#1;data_in = testData6[6300];
@(posedge clk);
#1;data_in = testData6[6301];
@(posedge clk);
#1;data_in = testData6[6302];
@(posedge clk);
#1;data_in = testData6[6303];
@(posedge clk);
#1;data_in = testData6[6304];
@(posedge clk);
#1;data_in = testData6[6305];
@(posedge clk);
#1;data_in = testData6[6306];
@(posedge clk);
#1;data_in = testData6[6307];
@(posedge clk);
#1;data_in = testData6[6308];
@(posedge clk);
#1;data_in = testData6[6309];
@(posedge clk);
#1;data_in = testData6[6310];
@(posedge clk);
#1;data_in = testData6[6311];
@(posedge clk);
#1;data_in = testData6[6312];
@(posedge clk);
#1;data_in = testData6[6313];
@(posedge clk);
#1;data_in = testData6[6314];
@(posedge clk);
#1;data_in = testData6[6315];
@(posedge clk);
#1;data_in = testData6[6316];
@(posedge clk);
#1;data_in = testData6[6317];
@(posedge clk);
#1;data_in = testData6[6318];
@(posedge clk);
#1;data_in = testData6[6319];
@(posedge clk);
#1;data_in = testData6[6320];
@(posedge clk);
#1;data_in = testData6[6321];
@(posedge clk);
#1;data_in = testData6[6322];
@(posedge clk);
#1;data_in = testData6[6323];
@(posedge clk);
#1;data_in = testData6[6324];
@(posedge clk);
#1;data_in = testData6[6325];
@(posedge clk);
#1;data_in = testData6[6326];
@(posedge clk);
#1;data_in = testData6[6327];
@(posedge clk);
#1;data_in = testData6[6328];
@(posedge clk);
#1;data_in = testData6[6329];
@(posedge clk);
#1;data_in = testData6[6330];
@(posedge clk);
#1;data_in = testData6[6331];
@(posedge clk);
#1;data_in = testData6[6332];
@(posedge clk);
#1;data_in = testData6[6333];
@(posedge clk);
#1;data_in = testData6[6334];
@(posedge clk);
#1;data_in = testData6[6335];
@(posedge clk);
#1;data_in = testData6[6336];
@(posedge clk);
#1;data_in = testData6[6337];
@(posedge clk);
#1;data_in = testData6[6338];
@(posedge clk);
#1;data_in = testData6[6339];
@(posedge clk);
#1;data_in = testData6[6340];
@(posedge clk);
#1;data_in = testData6[6341];
@(posedge clk);
#1;data_in = testData6[6342];
@(posedge clk);
#1;data_in = testData6[6343];
@(posedge clk);
#1;data_in = testData6[6344];
@(posedge clk);
#1;data_in = testData6[6345];
@(posedge clk);
#1;data_in = testData6[6346];
@(posedge clk);
#1;data_in = testData6[6347];
@(posedge clk);
#1;data_in = testData6[6348];
@(posedge clk);
#1;data_in = testData6[6349];
@(posedge clk);
#1;data_in = testData6[6350];
@(posedge clk);
#1;data_in = testData6[6351];
@(posedge clk);
#1;data_in = testData6[6352];
@(posedge clk);
#1;data_in = testData6[6353];
@(posedge clk);
#1;data_in = testData6[6354];
@(posedge clk);
#1;data_in = testData6[6355];
@(posedge clk);
#1;data_in = testData6[6356];
@(posedge clk);
#1;data_in = testData6[6357];
@(posedge clk);
#1;data_in = testData6[6358];
@(posedge clk);
#1;data_in = testData6[6359];
@(posedge clk);
#1;data_in = testData6[6360];
@(posedge clk);
#1;data_in = testData6[6361];
@(posedge clk);
#1;data_in = testData6[6362];
@(posedge clk);
#1;data_in = testData6[6363];
@(posedge clk);
#1;data_in = testData6[6364];
@(posedge clk);
#1;data_in = testData6[6365];
@(posedge clk);
#1;data_in = testData6[6366];
@(posedge clk);
#1;data_in = testData6[6367];
@(posedge clk);
#1;data_in = testData6[6368];
@(posedge clk);
#1;data_in = testData6[6369];
@(posedge clk);
#1;data_in = testData6[6370];
@(posedge clk);
#1;data_in = testData6[6371];
@(posedge clk);
#1;data_in = testData6[6372];
@(posedge clk);
#1;data_in = testData6[6373];
@(posedge clk);
#1;data_in = testData6[6374];
@(posedge clk);
#1;data_in = testData6[6375];
@(posedge clk);
#1;data_in = testData6[6376];
@(posedge clk);
#1;data_in = testData6[6377];
@(posedge clk);
#1;data_in = testData6[6378];
@(posedge clk);
#1;data_in = testData6[6379];
@(posedge clk);
#1;data_in = testData6[6380];
@(posedge clk);
#1;data_in = testData6[6381];
@(posedge clk);
#1;data_in = testData6[6382];
@(posedge clk);
#1;data_in = testData6[6383];
@(posedge clk);
#1;data_in = testData6[6384];
@(posedge clk);
#1;data_in = testData6[6385];
@(posedge clk);
#1;data_in = testData6[6386];
@(posedge clk);
#1;data_in = testData6[6387];
@(posedge clk);
#1;data_in = testData6[6388];
@(posedge clk);
#1;data_in = testData6[6389];
@(posedge clk);
#1;data_in = testData6[6390];
@(posedge clk);
#1;data_in = testData6[6391];
@(posedge clk);
#1;data_in = testData6[6392];
@(posedge clk);
#1;data_in = testData6[6393];
@(posedge clk);
#1;data_in = testData6[6394];
@(posedge clk);
#1;data_in = testData6[6395];
@(posedge clk);
#1;data_in = testData6[6396];
@(posedge clk);
#1;data_in = testData6[6397];
@(posedge clk);
#1;data_in = testData6[6398];
@(posedge clk);
#1;data_in = testData6[6399];
@(posedge clk);
#1;data_in = testData6[6400];
@(posedge clk);
#1;data_in = testData6[6401];
@(posedge clk);
#1;data_in = testData6[6402];
@(posedge clk);
#1;data_in = testData6[6403];
@(posedge clk);
#1;data_in = testData6[6404];
@(posedge clk);
#1;data_in = testData6[6405];
@(posedge clk);
#1;data_in = testData6[6406];
@(posedge clk);
#1;data_in = testData6[6407];
@(posedge clk);
#1;data_in = testData6[6408];
@(posedge clk);
#1;data_in = testData6[6409];
@(posedge clk);
#1;data_in = testData6[6410];
@(posedge clk);
#1;data_in = testData6[6411];
@(posedge clk);
#1;data_in = testData6[6412];
@(posedge clk);
#1;data_in = testData6[6413];
@(posedge clk);
#1;data_in = testData6[6414];
@(posedge clk);
#1;data_in = testData6[6415];
@(posedge clk);
#1;data_in = testData6[6416];
@(posedge clk);
#1;data_in = testData6[6417];
@(posedge clk);
#1;data_in = testData6[6418];
@(posedge clk);
#1;data_in = testData6[6419];
@(posedge clk);
#1;data_in = testData6[6420];
@(posedge clk);
#1;data_in = testData6[6421];
@(posedge clk);
#1;data_in = testData6[6422];
@(posedge clk);
#1;data_in = testData6[6423];
@(posedge clk);
#1;data_in = testData6[6424];
@(posedge clk);
#1;data_in = testData6[6425];
@(posedge clk);
#1;data_in = testData6[6426];
@(posedge clk);
#1;data_in = testData6[6427];
@(posedge clk);
#1;data_in = testData6[6428];
@(posedge clk);
#1;data_in = testData6[6429];
@(posedge clk);
#1;data_in = testData6[6430];
@(posedge clk);
#1;data_in = testData6[6431];
@(posedge clk);
#1;data_in = testData6[6432];
@(posedge clk);
#1;data_in = testData6[6433];
@(posedge clk);
#1;data_in = testData6[6434];
@(posedge clk);
#1;data_in = testData6[6435];
@(posedge clk);
#1;data_in = testData6[6436];
@(posedge clk);
#1;data_in = testData6[6437];
@(posedge clk);
#1;data_in = testData6[6438];
@(posedge clk);
#1;data_in = testData6[6439];
@(posedge clk);
#1;data_in = testData6[6440];
@(posedge clk);
#1;data_in = testData6[6441];
@(posedge clk);
#1;data_in = testData6[6442];
@(posedge clk);
#1;data_in = testData6[6443];
@(posedge clk);
#1;data_in = testData6[6444];
@(posedge clk);
#1;data_in = testData6[6445];
@(posedge clk);
#1;data_in = testData6[6446];
@(posedge clk);
#1;data_in = testData6[6447];
@(posedge clk);
#1;data_in = testData6[6448];
@(posedge clk);
#1;data_in = testData6[6449];
@(posedge clk);
#1;data_in = testData6[6450];
@(posedge clk);
#1;data_in = testData6[6451];
@(posedge clk);
#1;data_in = testData6[6452];
@(posedge clk);
#1;data_in = testData6[6453];
@(posedge clk);
#1;data_in = testData6[6454];
@(posedge clk);
#1;data_in = testData6[6455];
@(posedge clk);
#1;data_in = testData6[6456];
@(posedge clk);
#1;data_in = testData6[6457];
@(posedge clk);
#1;data_in = testData6[6458];
@(posedge clk);
#1;data_in = testData6[6459];
@(posedge clk);
#1;data_in = testData6[6460];
@(posedge clk);
#1;data_in = testData6[6461];
@(posedge clk);
#1;data_in = testData6[6462];
@(posedge clk);
#1;data_in = testData6[6463];
@(posedge clk);
#1;data_in = testData6[6464];
@(posedge clk);
#1;data_in = testData6[6465];
@(posedge clk);
#1;data_in = testData6[6466];
@(posedge clk);
#1;data_in = testData6[6467];
@(posedge clk);
#1;data_in = testData6[6468];
@(posedge clk);
#1;data_in = testData6[6469];
@(posedge clk);
#1;data_in = testData6[6470];
@(posedge clk);
#1;data_in = testData6[6471];
@(posedge clk);
#1;data_in = testData6[6472];
@(posedge clk);
#1;data_in = testData6[6473];
@(posedge clk);
#1;data_in = testData6[6474];
@(posedge clk);
#1;data_in = testData6[6475];
@(posedge clk);
#1;data_in = testData6[6476];
@(posedge clk);
#1;data_in = testData6[6477];
@(posedge clk);
#1;data_in = testData6[6478];
@(posedge clk);
#1;data_in = testData6[6479];
@(posedge clk);
#1;data_in = testData6[6480];
@(posedge clk);
#1;data_in = testData6[6481];
@(posedge clk);
#1;data_in = testData6[6482];
@(posedge clk);
#1;data_in = testData6[6483];
@(posedge clk);
#1;data_in = testData6[6484];
@(posedge clk);
#1;data_in = testData6[6485];
@(posedge clk);
#1;data_in = testData6[6486];
@(posedge clk);
#1;data_in = testData6[6487];
@(posedge clk);
#1;data_in = testData6[6488];
@(posedge clk);
#1;data_in = testData6[6489];
@(posedge clk);
#1;data_in = testData6[6490];
@(posedge clk);
#1;data_in = testData6[6491];
@(posedge clk);
#1;data_in = testData6[6492];
@(posedge clk);
#1;data_in = testData6[6493];
@(posedge clk);
#1;data_in = testData6[6494];
@(posedge clk);
#1;data_in = testData6[6495];
@(posedge clk);
#1;data_in = testData6[6496];
@(posedge clk);
#1;data_in = testData6[6497];
@(posedge clk);
#1;data_in = testData6[6498];
@(posedge clk);
#1;data_in = testData6[6499];
@(posedge clk);
#1;data_in = testData6[6500];
@(posedge clk);
#1;data_in = testData6[6501];
@(posedge clk);
#1;data_in = testData6[6502];
@(posedge clk);
#1;data_in = testData6[6503];
@(posedge clk);
#1;data_in = testData6[6504];
@(posedge clk);
#1;data_in = testData6[6505];
@(posedge clk);
#1;data_in = testData6[6506];
@(posedge clk);
#1;data_in = testData6[6507];
@(posedge clk);
#1;data_in = testData6[6508];
@(posedge clk);
#1;data_in = testData6[6509];
@(posedge clk);
#1;data_in = testData6[6510];
@(posedge clk);
#1;data_in = testData6[6511];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[6512]; 
@(posedge clk);
#1;data_in = testData6[6513];
@(posedge clk);
#1;data_in = testData6[6514];
@(posedge clk);
#1;data_in = testData6[6515];
@(posedge clk);
#1;data_in = testData6[6516];
@(posedge clk);
#1;data_in = testData6[6517];
@(posedge clk);
#1;data_in = testData6[6518];
@(posedge clk);
#1;data_in = testData6[6519];
@(posedge clk);
#1;data_in = testData6[6520];
@(posedge clk);
#1;data_in = testData6[6521];
@(posedge clk);
#1;data_in = testData6[6522];
@(posedge clk);
#1;data_in = testData6[6523];
@(posedge clk);
#1;data_in = testData6[6524];
@(posedge clk);
#1;data_in = testData6[6525];
@(posedge clk);
#1;data_in = testData6[6526];
@(posedge clk);
#1;data_in = testData6[6527];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[6528];
@(posedge clk);
#1;data_in = testData6[6529];
@(posedge clk);
#1;data_in = testData6[6530];
@(posedge clk);
#1;data_in = testData6[6531];
@(posedge clk);
#1;data_in = testData6[6532];
@(posedge clk);
#1;data_in = testData6[6533];
@(posedge clk);
#1;data_in = testData6[6534];
@(posedge clk);
#1;data_in = testData6[6535];
@(posedge clk);
#1;data_in = testData6[6536];
@(posedge clk);
#1;data_in = testData6[6537];
@(posedge clk);
#1;data_in = testData6[6538];
@(posedge clk);
#1;data_in = testData6[6539];
@(posedge clk);
#1;data_in = testData6[6540];
@(posedge clk);
#1;data_in = testData6[6541];
@(posedge clk);
#1;data_in = testData6[6542];
@(posedge clk);
#1;data_in = testData6[6543];
@(posedge clk);
#1;data_in = testData6[6544];
@(posedge clk);
#1;data_in = testData6[6545];
@(posedge clk);
#1;data_in = testData6[6546];
@(posedge clk);
#1;data_in = testData6[6547];
@(posedge clk);
#1;data_in = testData6[6548];
@(posedge clk);
#1;data_in = testData6[6549];
@(posedge clk);
#1;data_in = testData6[6550];
@(posedge clk);
#1;data_in = testData6[6551];
@(posedge clk);
#1;data_in = testData6[6552];
@(posedge clk);
#1;data_in = testData6[6553];
@(posedge clk);
#1;data_in = testData6[6554];
@(posedge clk);
#1;data_in = testData6[6555];
@(posedge clk);
#1;data_in = testData6[6556];
@(posedge clk);
#1;data_in = testData6[6557];
@(posedge clk);
#1;data_in = testData6[6558];
@(posedge clk);
#1;data_in = testData6[6559];
@(posedge clk);
#1;data_in = testData6[6560];
@(posedge clk);
#1;data_in = testData6[6561];
@(posedge clk);
#1;data_in = testData6[6562];
@(posedge clk);
#1;data_in = testData6[6563];
@(posedge clk);
#1;data_in = testData6[6564];
@(posedge clk);
#1;data_in = testData6[6565];
@(posedge clk);
#1;data_in = testData6[6566];
@(posedge clk);
#1;data_in = testData6[6567];
@(posedge clk);
#1;data_in = testData6[6568];
@(posedge clk);
#1;data_in = testData6[6569];
@(posedge clk);
#1;data_in = testData6[6570];
@(posedge clk);
#1;data_in = testData6[6571];
@(posedge clk);
#1;data_in = testData6[6572];
@(posedge clk);
#1;data_in = testData6[6573];
@(posedge clk);
#1;data_in = testData6[6574];
@(posedge clk);
#1;data_in = testData6[6575];
@(posedge clk);
#1;data_in = testData6[6576];
@(posedge clk);
#1;data_in = testData6[6577];
@(posedge clk);
#1;data_in = testData6[6578];
@(posedge clk);
#1;data_in = testData6[6579];
@(posedge clk);
#1;data_in = testData6[6580];
@(posedge clk);
#1;data_in = testData6[6581];
@(posedge clk);
#1;data_in = testData6[6582];
@(posedge clk);
#1;data_in = testData6[6583];
@(posedge clk);
#1;data_in = testData6[6584];
@(posedge clk);
#1;data_in = testData6[6585];
@(posedge clk);
#1;data_in = testData6[6586];
@(posedge clk);
#1;data_in = testData6[6587];
@(posedge clk);
#1;data_in = testData6[6588];
@(posedge clk);
#1;data_in = testData6[6589];
@(posedge clk);
#1;data_in = testData6[6590];
@(posedge clk);
#1;data_in = testData6[6591];
@(posedge clk);
#1;data_in = testData6[6592];
@(posedge clk);
#1;data_in = testData6[6593];
@(posedge clk);
#1;data_in = testData6[6594];
@(posedge clk);
#1;data_in = testData6[6595];
@(posedge clk);
#1;data_in = testData6[6596];
@(posedge clk);
#1;data_in = testData6[6597];
@(posedge clk);
#1;data_in = testData6[6598];
@(posedge clk);
#1;data_in = testData6[6599];
@(posedge clk);
#1;data_in = testData6[6600];
@(posedge clk);
#1;data_in = testData6[6601];
@(posedge clk);
#1;data_in = testData6[6602];
@(posedge clk);
#1;data_in = testData6[6603];
@(posedge clk);
#1;data_in = testData6[6604];
@(posedge clk);
#1;data_in = testData6[6605];
@(posedge clk);
#1;data_in = testData6[6606];
@(posedge clk);
#1;data_in = testData6[6607];
@(posedge clk);
#1;data_in = testData6[6608];
@(posedge clk);
#1;data_in = testData6[6609];
@(posedge clk);
#1;data_in = testData6[6610];
@(posedge clk);
#1;data_in = testData6[6611];
@(posedge clk);
#1;data_in = testData6[6612];
@(posedge clk);
#1;data_in = testData6[6613];
@(posedge clk);
#1;data_in = testData6[6614];
@(posedge clk);
#1;data_in = testData6[6615];
@(posedge clk);
#1;data_in = testData6[6616];
@(posedge clk);
#1;data_in = testData6[6617];
@(posedge clk);
#1;data_in = testData6[6618];
@(posedge clk);
#1;data_in = testData6[6619];
@(posedge clk);
#1;data_in = testData6[6620];
@(posedge clk);
#1;data_in = testData6[6621];
@(posedge clk);
#1;data_in = testData6[6622];
@(posedge clk);
#1;data_in = testData6[6623];
@(posedge clk);
#1;data_in = testData6[6624];
@(posedge clk);
#1;data_in = testData6[6625];
@(posedge clk);
#1;data_in = testData6[6626];
@(posedge clk);
#1;data_in = testData6[6627];
@(posedge clk);
#1;data_in = testData6[6628];
@(posedge clk);
#1;data_in = testData6[6629];
@(posedge clk);
#1;data_in = testData6[6630];
@(posedge clk);
#1;data_in = testData6[6631];
@(posedge clk);
#1;data_in = testData6[6632];
@(posedge clk);
#1;data_in = testData6[6633];
@(posedge clk);
#1;data_in = testData6[6634];
@(posedge clk);
#1;data_in = testData6[6635];
@(posedge clk);
#1;data_in = testData6[6636];
@(posedge clk);
#1;data_in = testData6[6637];
@(posedge clk);
#1;data_in = testData6[6638];
@(posedge clk);
#1;data_in = testData6[6639];
@(posedge clk);
#1;data_in = testData6[6640];
@(posedge clk);
#1;data_in = testData6[6641];
@(posedge clk);
#1;data_in = testData6[6642];
@(posedge clk);
#1;data_in = testData6[6643];
@(posedge clk);
#1;data_in = testData6[6644];
@(posedge clk);
#1;data_in = testData6[6645];
@(posedge clk);
#1;data_in = testData6[6646];
@(posedge clk);
#1;data_in = testData6[6647];
@(posedge clk);
#1;data_in = testData6[6648];
@(posedge clk);
#1;data_in = testData6[6649];
@(posedge clk);
#1;data_in = testData6[6650];
@(posedge clk);
#1;data_in = testData6[6651];
@(posedge clk);
#1;data_in = testData6[6652];
@(posedge clk);
#1;data_in = testData6[6653];
@(posedge clk);
#1;data_in = testData6[6654];
@(posedge clk);
#1;data_in = testData6[6655];
@(posedge clk);
#1;data_in = testData6[6656];
@(posedge clk);
#1;data_in = testData6[6657];
@(posedge clk);
#1;data_in = testData6[6658];
@(posedge clk);
#1;data_in = testData6[6659];
@(posedge clk);
#1;data_in = testData6[6660];
@(posedge clk);
#1;data_in = testData6[6661];
@(posedge clk);
#1;data_in = testData6[6662];
@(posedge clk);
#1;data_in = testData6[6663];
@(posedge clk);
#1;data_in = testData6[6664];
@(posedge clk);
#1;data_in = testData6[6665];
@(posedge clk);
#1;data_in = testData6[6666];
@(posedge clk);
#1;data_in = testData6[6667];
@(posedge clk);
#1;data_in = testData6[6668];
@(posedge clk);
#1;data_in = testData6[6669];
@(posedge clk);
#1;data_in = testData6[6670];
@(posedge clk);
#1;data_in = testData6[6671];
@(posedge clk);
#1;data_in = testData6[6672];
@(posedge clk);
#1;data_in = testData6[6673];
@(posedge clk);
#1;data_in = testData6[6674];
@(posedge clk);
#1;data_in = testData6[6675];
@(posedge clk);
#1;data_in = testData6[6676];
@(posedge clk);
#1;data_in = testData6[6677];
@(posedge clk);
#1;data_in = testData6[6678];
@(posedge clk);
#1;data_in = testData6[6679];
@(posedge clk);
#1;data_in = testData6[6680];
@(posedge clk);
#1;data_in = testData6[6681];
@(posedge clk);
#1;data_in = testData6[6682];
@(posedge clk);
#1;data_in = testData6[6683];
@(posedge clk);
#1;data_in = testData6[6684];
@(posedge clk);
#1;data_in = testData6[6685];
@(posedge clk);
#1;data_in = testData6[6686];
@(posedge clk);
#1;data_in = testData6[6687];
@(posedge clk);
#1;data_in = testData6[6688];
@(posedge clk);
#1;data_in = testData6[6689];
@(posedge clk);
#1;data_in = testData6[6690];
@(posedge clk);
#1;data_in = testData6[6691];
@(posedge clk);
#1;data_in = testData6[6692];
@(posedge clk);
#1;data_in = testData6[6693];
@(posedge clk);
#1;data_in = testData6[6694];
@(posedge clk);
#1;data_in = testData6[6695];
@(posedge clk);
#1;data_in = testData6[6696];
@(posedge clk);
#1;data_in = testData6[6697];
@(posedge clk);
#1;data_in = testData6[6698];
@(posedge clk);
#1;data_in = testData6[6699];
@(posedge clk);
#1;data_in = testData6[6700];
@(posedge clk);
#1;data_in = testData6[6701];
@(posedge clk);
#1;data_in = testData6[6702];
@(posedge clk);
#1;data_in = testData6[6703];
@(posedge clk);
#1;data_in = testData6[6704];
@(posedge clk);
#1;data_in = testData6[6705];
@(posedge clk);
#1;data_in = testData6[6706];
@(posedge clk);
#1;data_in = testData6[6707];
@(posedge clk);
#1;data_in = testData6[6708];
@(posedge clk);
#1;data_in = testData6[6709];
@(posedge clk);
#1;data_in = testData6[6710];
@(posedge clk);
#1;data_in = testData6[6711];
@(posedge clk);
#1;data_in = testData6[6712];
@(posedge clk);
#1;data_in = testData6[6713];
@(posedge clk);
#1;data_in = testData6[6714];
@(posedge clk);
#1;data_in = testData6[6715];
@(posedge clk);
#1;data_in = testData6[6716];
@(posedge clk);
#1;data_in = testData6[6717];
@(posedge clk);
#1;data_in = testData6[6718];
@(posedge clk);
#1;data_in = testData6[6719];
@(posedge clk);
#1;data_in = testData6[6720];
@(posedge clk);
#1;data_in = testData6[6721];
@(posedge clk);
#1;data_in = testData6[6722];
@(posedge clk);
#1;data_in = testData6[6723];
@(posedge clk);
#1;data_in = testData6[6724];
@(posedge clk);
#1;data_in = testData6[6725];
@(posedge clk);
#1;data_in = testData6[6726];
@(posedge clk);
#1;data_in = testData6[6727];
@(posedge clk);
#1;data_in = testData6[6728];
@(posedge clk);
#1;data_in = testData6[6729];
@(posedge clk);
#1;data_in = testData6[6730];
@(posedge clk);
#1;data_in = testData6[6731];
@(posedge clk);
#1;data_in = testData6[6732];
@(posedge clk);
#1;data_in = testData6[6733];
@(posedge clk);
#1;data_in = testData6[6734];
@(posedge clk);
#1;data_in = testData6[6735];
@(posedge clk);
#1;data_in = testData6[6736];
@(posedge clk);
#1;data_in = testData6[6737];
@(posedge clk);
#1;data_in = testData6[6738];
@(posedge clk);
#1;data_in = testData6[6739];
@(posedge clk);
#1;data_in = testData6[6740];
@(posedge clk);
#1;data_in = testData6[6741];
@(posedge clk);
#1;data_in = testData6[6742];
@(posedge clk);
#1;data_in = testData6[6743];
@(posedge clk);
#1;data_in = testData6[6744];
@(posedge clk);
#1;data_in = testData6[6745];
@(posedge clk);
#1;data_in = testData6[6746];
@(posedge clk);
#1;data_in = testData6[6747];
@(posedge clk);
#1;data_in = testData6[6748];
@(posedge clk);
#1;data_in = testData6[6749];
@(posedge clk);
#1;data_in = testData6[6750];
@(posedge clk);
#1;data_in = testData6[6751];
@(posedge clk);
#1;data_in = testData6[6752];
@(posedge clk);
#1;data_in = testData6[6753];
@(posedge clk);
#1;data_in = testData6[6754];
@(posedge clk);
#1;data_in = testData6[6755];
@(posedge clk);
#1;data_in = testData6[6756];
@(posedge clk);
#1;data_in = testData6[6757];
@(posedge clk);
#1;data_in = testData6[6758];
@(posedge clk);
#1;data_in = testData6[6759];
@(posedge clk);
#1;data_in = testData6[6760];
@(posedge clk);
#1;data_in = testData6[6761];
@(posedge clk);
#1;data_in = testData6[6762];
@(posedge clk);
#1;data_in = testData6[6763];
@(posedge clk);
#1;data_in = testData6[6764];
@(posedge clk);
#1;data_in = testData6[6765];
@(posedge clk);
#1;data_in = testData6[6766];
@(posedge clk);
#1;data_in = testData6[6767];
@(posedge clk);
#1;data_in = testData6[6768];
@(posedge clk);
#1;data_in = testData6[6769];
@(posedge clk);
#1;data_in = testData6[6770];
@(posedge clk);
#1;data_in = testData6[6771];
@(posedge clk);
#1;data_in = testData6[6772];
@(posedge clk);
#1;data_in = testData6[6773];
@(posedge clk);
#1;data_in = testData6[6774];
@(posedge clk);
#1;data_in = testData6[6775];
@(posedge clk);
#1;data_in = testData6[6776];
@(posedge clk);
#1;data_in = testData6[6777];
@(posedge clk);
#1;data_in = testData6[6778];
@(posedge clk);
#1;data_in = testData6[6779];
@(posedge clk);
#1;data_in = testData6[6780];
@(posedge clk);
#1;data_in = testData6[6781];
@(posedge clk);
#1;data_in = testData6[6782];
@(posedge clk);
#1;data_in = testData6[6783];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[6784]; 
@(posedge clk);
#1;data_in = testData6[6785];
@(posedge clk);
#1;data_in = testData6[6786];
@(posedge clk);
#1;data_in = testData6[6787];
@(posedge clk);
#1;data_in = testData6[6788];
@(posedge clk);
#1;data_in = testData6[6789];
@(posedge clk);
#1;data_in = testData6[6790];
@(posedge clk);
#1;data_in = testData6[6791];
@(posedge clk);
#1;data_in = testData6[6792];
@(posedge clk);
#1;data_in = testData6[6793];
@(posedge clk);
#1;data_in = testData6[6794];
@(posedge clk);
#1;data_in = testData6[6795];
@(posedge clk);
#1;data_in = testData6[6796];
@(posedge clk);
#1;data_in = testData6[6797];
@(posedge clk);
#1;data_in = testData6[6798];
@(posedge clk);
#1;data_in = testData6[6799];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[6800];
@(posedge clk);
#1;data_in = testData6[6801];
@(posedge clk);
#1;data_in = testData6[6802];
@(posedge clk);
#1;data_in = testData6[6803];
@(posedge clk);
#1;data_in = testData6[6804];
@(posedge clk);
#1;data_in = testData6[6805];
@(posedge clk);
#1;data_in = testData6[6806];
@(posedge clk);
#1;data_in = testData6[6807];
@(posedge clk);
#1;data_in = testData6[6808];
@(posedge clk);
#1;data_in = testData6[6809];
@(posedge clk);
#1;data_in = testData6[6810];
@(posedge clk);
#1;data_in = testData6[6811];
@(posedge clk);
#1;data_in = testData6[6812];
@(posedge clk);
#1;data_in = testData6[6813];
@(posedge clk);
#1;data_in = testData6[6814];
@(posedge clk);
#1;data_in = testData6[6815];
@(posedge clk);
#1;data_in = testData6[6816];
@(posedge clk);
#1;data_in = testData6[6817];
@(posedge clk);
#1;data_in = testData6[6818];
@(posedge clk);
#1;data_in = testData6[6819];
@(posedge clk);
#1;data_in = testData6[6820];
@(posedge clk);
#1;data_in = testData6[6821];
@(posedge clk);
#1;data_in = testData6[6822];
@(posedge clk);
#1;data_in = testData6[6823];
@(posedge clk);
#1;data_in = testData6[6824];
@(posedge clk);
#1;data_in = testData6[6825];
@(posedge clk);
#1;data_in = testData6[6826];
@(posedge clk);
#1;data_in = testData6[6827];
@(posedge clk);
#1;data_in = testData6[6828];
@(posedge clk);
#1;data_in = testData6[6829];
@(posedge clk);
#1;data_in = testData6[6830];
@(posedge clk);
#1;data_in = testData6[6831];
@(posedge clk);
#1;data_in = testData6[6832];
@(posedge clk);
#1;data_in = testData6[6833];
@(posedge clk);
#1;data_in = testData6[6834];
@(posedge clk);
#1;data_in = testData6[6835];
@(posedge clk);
#1;data_in = testData6[6836];
@(posedge clk);
#1;data_in = testData6[6837];
@(posedge clk);
#1;data_in = testData6[6838];
@(posedge clk);
#1;data_in = testData6[6839];
@(posedge clk);
#1;data_in = testData6[6840];
@(posedge clk);
#1;data_in = testData6[6841];
@(posedge clk);
#1;data_in = testData6[6842];
@(posedge clk);
#1;data_in = testData6[6843];
@(posedge clk);
#1;data_in = testData6[6844];
@(posedge clk);
#1;data_in = testData6[6845];
@(posedge clk);
#1;data_in = testData6[6846];
@(posedge clk);
#1;data_in = testData6[6847];
@(posedge clk);
#1;data_in = testData6[6848];
@(posedge clk);
#1;data_in = testData6[6849];
@(posedge clk);
#1;data_in = testData6[6850];
@(posedge clk);
#1;data_in = testData6[6851];
@(posedge clk);
#1;data_in = testData6[6852];
@(posedge clk);
#1;data_in = testData6[6853];
@(posedge clk);
#1;data_in = testData6[6854];
@(posedge clk);
#1;data_in = testData6[6855];
@(posedge clk);
#1;data_in = testData6[6856];
@(posedge clk);
#1;data_in = testData6[6857];
@(posedge clk);
#1;data_in = testData6[6858];
@(posedge clk);
#1;data_in = testData6[6859];
@(posedge clk);
#1;data_in = testData6[6860];
@(posedge clk);
#1;data_in = testData6[6861];
@(posedge clk);
#1;data_in = testData6[6862];
@(posedge clk);
#1;data_in = testData6[6863];
@(posedge clk);
#1;data_in = testData6[6864];
@(posedge clk);
#1;data_in = testData6[6865];
@(posedge clk);
#1;data_in = testData6[6866];
@(posedge clk);
#1;data_in = testData6[6867];
@(posedge clk);
#1;data_in = testData6[6868];
@(posedge clk);
#1;data_in = testData6[6869];
@(posedge clk);
#1;data_in = testData6[6870];
@(posedge clk);
#1;data_in = testData6[6871];
@(posedge clk);
#1;data_in = testData6[6872];
@(posedge clk);
#1;data_in = testData6[6873];
@(posedge clk);
#1;data_in = testData6[6874];
@(posedge clk);
#1;data_in = testData6[6875];
@(posedge clk);
#1;data_in = testData6[6876];
@(posedge clk);
#1;data_in = testData6[6877];
@(posedge clk);
#1;data_in = testData6[6878];
@(posedge clk);
#1;data_in = testData6[6879];
@(posedge clk);
#1;data_in = testData6[6880];
@(posedge clk);
#1;data_in = testData6[6881];
@(posedge clk);
#1;data_in = testData6[6882];
@(posedge clk);
#1;data_in = testData6[6883];
@(posedge clk);
#1;data_in = testData6[6884];
@(posedge clk);
#1;data_in = testData6[6885];
@(posedge clk);
#1;data_in = testData6[6886];
@(posedge clk);
#1;data_in = testData6[6887];
@(posedge clk);
#1;data_in = testData6[6888];
@(posedge clk);
#1;data_in = testData6[6889];
@(posedge clk);
#1;data_in = testData6[6890];
@(posedge clk);
#1;data_in = testData6[6891];
@(posedge clk);
#1;data_in = testData6[6892];
@(posedge clk);
#1;data_in = testData6[6893];
@(posedge clk);
#1;data_in = testData6[6894];
@(posedge clk);
#1;data_in = testData6[6895];
@(posedge clk);
#1;data_in = testData6[6896];
@(posedge clk);
#1;data_in = testData6[6897];
@(posedge clk);
#1;data_in = testData6[6898];
@(posedge clk);
#1;data_in = testData6[6899];
@(posedge clk);
#1;data_in = testData6[6900];
@(posedge clk);
#1;data_in = testData6[6901];
@(posedge clk);
#1;data_in = testData6[6902];
@(posedge clk);
#1;data_in = testData6[6903];
@(posedge clk);
#1;data_in = testData6[6904];
@(posedge clk);
#1;data_in = testData6[6905];
@(posedge clk);
#1;data_in = testData6[6906];
@(posedge clk);
#1;data_in = testData6[6907];
@(posedge clk);
#1;data_in = testData6[6908];
@(posedge clk);
#1;data_in = testData6[6909];
@(posedge clk);
#1;data_in = testData6[6910];
@(posedge clk);
#1;data_in = testData6[6911];
@(posedge clk);
#1;data_in = testData6[6912];
@(posedge clk);
#1;data_in = testData6[6913];
@(posedge clk);
#1;data_in = testData6[6914];
@(posedge clk);
#1;data_in = testData6[6915];
@(posedge clk);
#1;data_in = testData6[6916];
@(posedge clk);
#1;data_in = testData6[6917];
@(posedge clk);
#1;data_in = testData6[6918];
@(posedge clk);
#1;data_in = testData6[6919];
@(posedge clk);
#1;data_in = testData6[6920];
@(posedge clk);
#1;data_in = testData6[6921];
@(posedge clk);
#1;data_in = testData6[6922];
@(posedge clk);
#1;data_in = testData6[6923];
@(posedge clk);
#1;data_in = testData6[6924];
@(posedge clk);
#1;data_in = testData6[6925];
@(posedge clk);
#1;data_in = testData6[6926];
@(posedge clk);
#1;data_in = testData6[6927];
@(posedge clk);
#1;data_in = testData6[6928];
@(posedge clk);
#1;data_in = testData6[6929];
@(posedge clk);
#1;data_in = testData6[6930];
@(posedge clk);
#1;data_in = testData6[6931];
@(posedge clk);
#1;data_in = testData6[6932];
@(posedge clk);
#1;data_in = testData6[6933];
@(posedge clk);
#1;data_in = testData6[6934];
@(posedge clk);
#1;data_in = testData6[6935];
@(posedge clk);
#1;data_in = testData6[6936];
@(posedge clk);
#1;data_in = testData6[6937];
@(posedge clk);
#1;data_in = testData6[6938];
@(posedge clk);
#1;data_in = testData6[6939];
@(posedge clk);
#1;data_in = testData6[6940];
@(posedge clk);
#1;data_in = testData6[6941];
@(posedge clk);
#1;data_in = testData6[6942];
@(posedge clk);
#1;data_in = testData6[6943];
@(posedge clk);
#1;data_in = testData6[6944];
@(posedge clk);
#1;data_in = testData6[6945];
@(posedge clk);
#1;data_in = testData6[6946];
@(posedge clk);
#1;data_in = testData6[6947];
@(posedge clk);
#1;data_in = testData6[6948];
@(posedge clk);
#1;data_in = testData6[6949];
@(posedge clk);
#1;data_in = testData6[6950];
@(posedge clk);
#1;data_in = testData6[6951];
@(posedge clk);
#1;data_in = testData6[6952];
@(posedge clk);
#1;data_in = testData6[6953];
@(posedge clk);
#1;data_in = testData6[6954];
@(posedge clk);
#1;data_in = testData6[6955];
@(posedge clk);
#1;data_in = testData6[6956];
@(posedge clk);
#1;data_in = testData6[6957];
@(posedge clk);
#1;data_in = testData6[6958];
@(posedge clk);
#1;data_in = testData6[6959];
@(posedge clk);
#1;data_in = testData6[6960];
@(posedge clk);
#1;data_in = testData6[6961];
@(posedge clk);
#1;data_in = testData6[6962];
@(posedge clk);
#1;data_in = testData6[6963];
@(posedge clk);
#1;data_in = testData6[6964];
@(posedge clk);
#1;data_in = testData6[6965];
@(posedge clk);
#1;data_in = testData6[6966];
@(posedge clk);
#1;data_in = testData6[6967];
@(posedge clk);
#1;data_in = testData6[6968];
@(posedge clk);
#1;data_in = testData6[6969];
@(posedge clk);
#1;data_in = testData6[6970];
@(posedge clk);
#1;data_in = testData6[6971];
@(posedge clk);
#1;data_in = testData6[6972];
@(posedge clk);
#1;data_in = testData6[6973];
@(posedge clk);
#1;data_in = testData6[6974];
@(posedge clk);
#1;data_in = testData6[6975];
@(posedge clk);
#1;data_in = testData6[6976];
@(posedge clk);
#1;data_in = testData6[6977];
@(posedge clk);
#1;data_in = testData6[6978];
@(posedge clk);
#1;data_in = testData6[6979];
@(posedge clk);
#1;data_in = testData6[6980];
@(posedge clk);
#1;data_in = testData6[6981];
@(posedge clk);
#1;data_in = testData6[6982];
@(posedge clk);
#1;data_in = testData6[6983];
@(posedge clk);
#1;data_in = testData6[6984];
@(posedge clk);
#1;data_in = testData6[6985];
@(posedge clk);
#1;data_in = testData6[6986];
@(posedge clk);
#1;data_in = testData6[6987];
@(posedge clk);
#1;data_in = testData6[6988];
@(posedge clk);
#1;data_in = testData6[6989];
@(posedge clk);
#1;data_in = testData6[6990];
@(posedge clk);
#1;data_in = testData6[6991];
@(posedge clk);
#1;data_in = testData6[6992];
@(posedge clk);
#1;data_in = testData6[6993];
@(posedge clk);
#1;data_in = testData6[6994];
@(posedge clk);
#1;data_in = testData6[6995];
@(posedge clk);
#1;data_in = testData6[6996];
@(posedge clk);
#1;data_in = testData6[6997];
@(posedge clk);
#1;data_in = testData6[6998];
@(posedge clk);
#1;data_in = testData6[6999];
@(posedge clk);
#1;data_in = testData6[7000];
@(posedge clk);
#1;data_in = testData6[7001];
@(posedge clk);
#1;data_in = testData6[7002];
@(posedge clk);
#1;data_in = testData6[7003];
@(posedge clk);
#1;data_in = testData6[7004];
@(posedge clk);
#1;data_in = testData6[7005];
@(posedge clk);
#1;data_in = testData6[7006];
@(posedge clk);
#1;data_in = testData6[7007];
@(posedge clk);
#1;data_in = testData6[7008];
@(posedge clk);
#1;data_in = testData6[7009];
@(posedge clk);
#1;data_in = testData6[7010];
@(posedge clk);
#1;data_in = testData6[7011];
@(posedge clk);
#1;data_in = testData6[7012];
@(posedge clk);
#1;data_in = testData6[7013];
@(posedge clk);
#1;data_in = testData6[7014];
@(posedge clk);
#1;data_in = testData6[7015];
@(posedge clk);
#1;data_in = testData6[7016];
@(posedge clk);
#1;data_in = testData6[7017];
@(posedge clk);
#1;data_in = testData6[7018];
@(posedge clk);
#1;data_in = testData6[7019];
@(posedge clk);
#1;data_in = testData6[7020];
@(posedge clk);
#1;data_in = testData6[7021];
@(posedge clk);
#1;data_in = testData6[7022];
@(posedge clk);
#1;data_in = testData6[7023];
@(posedge clk);
#1;data_in = testData6[7024];
@(posedge clk);
#1;data_in = testData6[7025];
@(posedge clk);
#1;data_in = testData6[7026];
@(posedge clk);
#1;data_in = testData6[7027];
@(posedge clk);
#1;data_in = testData6[7028];
@(posedge clk);
#1;data_in = testData6[7029];
@(posedge clk);
#1;data_in = testData6[7030];
@(posedge clk);
#1;data_in = testData6[7031];
@(posedge clk);
#1;data_in = testData6[7032];
@(posedge clk);
#1;data_in = testData6[7033];
@(posedge clk);
#1;data_in = testData6[7034];
@(posedge clk);
#1;data_in = testData6[7035];
@(posedge clk);
#1;data_in = testData6[7036];
@(posedge clk);
#1;data_in = testData6[7037];
@(posedge clk);
#1;data_in = testData6[7038];
@(posedge clk);
#1;data_in = testData6[7039];
@(posedge clk);
#1;data_in = testData6[7040];
@(posedge clk);
#1;data_in = testData6[7041];
@(posedge clk);
#1;data_in = testData6[7042];
@(posedge clk);
#1;data_in = testData6[7043];
@(posedge clk);
#1;data_in = testData6[7044];
@(posedge clk);
#1;data_in = testData6[7045];
@(posedge clk);
#1;data_in = testData6[7046];
@(posedge clk);
#1;data_in = testData6[7047];
@(posedge clk);
#1;data_in = testData6[7048];
@(posedge clk);
#1;data_in = testData6[7049];
@(posedge clk);
#1;data_in = testData6[7050];
@(posedge clk);
#1;data_in = testData6[7051];
@(posedge clk);
#1;data_in = testData6[7052];
@(posedge clk);
#1;data_in = testData6[7053];
@(posedge clk);
#1;data_in = testData6[7054];
@(posedge clk);
#1;data_in = testData6[7055];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[7056]; 
@(posedge clk);
#1;data_in = testData6[7057];
@(posedge clk);
#1;data_in = testData6[7058];
@(posedge clk);
#1;data_in = testData6[7059];
@(posedge clk);
#1;data_in = testData6[7060];
@(posedge clk);
#1;data_in = testData6[7061];
@(posedge clk);
#1;data_in = testData6[7062];
@(posedge clk);
#1;data_in = testData6[7063];
@(posedge clk);
#1;data_in = testData6[7064];
@(posedge clk);
#1;data_in = testData6[7065];
@(posedge clk);
#1;data_in = testData6[7066];
@(posedge clk);
#1;data_in = testData6[7067];
@(posedge clk);
#1;data_in = testData6[7068];
@(posedge clk);
#1;data_in = testData6[7069];
@(posedge clk);
#1;data_in = testData6[7070];
@(posedge clk);
#1;data_in = testData6[7071];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[7072];
@(posedge clk);
#1;data_in = testData6[7073];
@(posedge clk);
#1;data_in = testData6[7074];
@(posedge clk);
#1;data_in = testData6[7075];
@(posedge clk);
#1;data_in = testData6[7076];
@(posedge clk);
#1;data_in = testData6[7077];
@(posedge clk);
#1;data_in = testData6[7078];
@(posedge clk);
#1;data_in = testData6[7079];
@(posedge clk);
#1;data_in = testData6[7080];
@(posedge clk);
#1;data_in = testData6[7081];
@(posedge clk);
#1;data_in = testData6[7082];
@(posedge clk);
#1;data_in = testData6[7083];
@(posedge clk);
#1;data_in = testData6[7084];
@(posedge clk);
#1;data_in = testData6[7085];
@(posedge clk);
#1;data_in = testData6[7086];
@(posedge clk);
#1;data_in = testData6[7087];
@(posedge clk);
#1;data_in = testData6[7088];
@(posedge clk);
#1;data_in = testData6[7089];
@(posedge clk);
#1;data_in = testData6[7090];
@(posedge clk);
#1;data_in = testData6[7091];
@(posedge clk);
#1;data_in = testData6[7092];
@(posedge clk);
#1;data_in = testData6[7093];
@(posedge clk);
#1;data_in = testData6[7094];
@(posedge clk);
#1;data_in = testData6[7095];
@(posedge clk);
#1;data_in = testData6[7096];
@(posedge clk);
#1;data_in = testData6[7097];
@(posedge clk);
#1;data_in = testData6[7098];
@(posedge clk);
#1;data_in = testData6[7099];
@(posedge clk);
#1;data_in = testData6[7100];
@(posedge clk);
#1;data_in = testData6[7101];
@(posedge clk);
#1;data_in = testData6[7102];
@(posedge clk);
#1;data_in = testData6[7103];
@(posedge clk);
#1;data_in = testData6[7104];
@(posedge clk);
#1;data_in = testData6[7105];
@(posedge clk);
#1;data_in = testData6[7106];
@(posedge clk);
#1;data_in = testData6[7107];
@(posedge clk);
#1;data_in = testData6[7108];
@(posedge clk);
#1;data_in = testData6[7109];
@(posedge clk);
#1;data_in = testData6[7110];
@(posedge clk);
#1;data_in = testData6[7111];
@(posedge clk);
#1;data_in = testData6[7112];
@(posedge clk);
#1;data_in = testData6[7113];
@(posedge clk);
#1;data_in = testData6[7114];
@(posedge clk);
#1;data_in = testData6[7115];
@(posedge clk);
#1;data_in = testData6[7116];
@(posedge clk);
#1;data_in = testData6[7117];
@(posedge clk);
#1;data_in = testData6[7118];
@(posedge clk);
#1;data_in = testData6[7119];
@(posedge clk);
#1;data_in = testData6[7120];
@(posedge clk);
#1;data_in = testData6[7121];
@(posedge clk);
#1;data_in = testData6[7122];
@(posedge clk);
#1;data_in = testData6[7123];
@(posedge clk);
#1;data_in = testData6[7124];
@(posedge clk);
#1;data_in = testData6[7125];
@(posedge clk);
#1;data_in = testData6[7126];
@(posedge clk);
#1;data_in = testData6[7127];
@(posedge clk);
#1;data_in = testData6[7128];
@(posedge clk);
#1;data_in = testData6[7129];
@(posedge clk);
#1;data_in = testData6[7130];
@(posedge clk);
#1;data_in = testData6[7131];
@(posedge clk);
#1;data_in = testData6[7132];
@(posedge clk);
#1;data_in = testData6[7133];
@(posedge clk);
#1;data_in = testData6[7134];
@(posedge clk);
#1;data_in = testData6[7135];
@(posedge clk);
#1;data_in = testData6[7136];
@(posedge clk);
#1;data_in = testData6[7137];
@(posedge clk);
#1;data_in = testData6[7138];
@(posedge clk);
#1;data_in = testData6[7139];
@(posedge clk);
#1;data_in = testData6[7140];
@(posedge clk);
#1;data_in = testData6[7141];
@(posedge clk);
#1;data_in = testData6[7142];
@(posedge clk);
#1;data_in = testData6[7143];
@(posedge clk);
#1;data_in = testData6[7144];
@(posedge clk);
#1;data_in = testData6[7145];
@(posedge clk);
#1;data_in = testData6[7146];
@(posedge clk);
#1;data_in = testData6[7147];
@(posedge clk);
#1;data_in = testData6[7148];
@(posedge clk);
#1;data_in = testData6[7149];
@(posedge clk);
#1;data_in = testData6[7150];
@(posedge clk);
#1;data_in = testData6[7151];
@(posedge clk);
#1;data_in = testData6[7152];
@(posedge clk);
#1;data_in = testData6[7153];
@(posedge clk);
#1;data_in = testData6[7154];
@(posedge clk);
#1;data_in = testData6[7155];
@(posedge clk);
#1;data_in = testData6[7156];
@(posedge clk);
#1;data_in = testData6[7157];
@(posedge clk);
#1;data_in = testData6[7158];
@(posedge clk);
#1;data_in = testData6[7159];
@(posedge clk);
#1;data_in = testData6[7160];
@(posedge clk);
#1;data_in = testData6[7161];
@(posedge clk);
#1;data_in = testData6[7162];
@(posedge clk);
#1;data_in = testData6[7163];
@(posedge clk);
#1;data_in = testData6[7164];
@(posedge clk);
#1;data_in = testData6[7165];
@(posedge clk);
#1;data_in = testData6[7166];
@(posedge clk);
#1;data_in = testData6[7167];
@(posedge clk);
#1;data_in = testData6[7168];
@(posedge clk);
#1;data_in = testData6[7169];
@(posedge clk);
#1;data_in = testData6[7170];
@(posedge clk);
#1;data_in = testData6[7171];
@(posedge clk);
#1;data_in = testData6[7172];
@(posedge clk);
#1;data_in = testData6[7173];
@(posedge clk);
#1;data_in = testData6[7174];
@(posedge clk);
#1;data_in = testData6[7175];
@(posedge clk);
#1;data_in = testData6[7176];
@(posedge clk);
#1;data_in = testData6[7177];
@(posedge clk);
#1;data_in = testData6[7178];
@(posedge clk);
#1;data_in = testData6[7179];
@(posedge clk);
#1;data_in = testData6[7180];
@(posedge clk);
#1;data_in = testData6[7181];
@(posedge clk);
#1;data_in = testData6[7182];
@(posedge clk);
#1;data_in = testData6[7183];
@(posedge clk);
#1;data_in = testData6[7184];
@(posedge clk);
#1;data_in = testData6[7185];
@(posedge clk);
#1;data_in = testData6[7186];
@(posedge clk);
#1;data_in = testData6[7187];
@(posedge clk);
#1;data_in = testData6[7188];
@(posedge clk);
#1;data_in = testData6[7189];
@(posedge clk);
#1;data_in = testData6[7190];
@(posedge clk);
#1;data_in = testData6[7191];
@(posedge clk);
#1;data_in = testData6[7192];
@(posedge clk);
#1;data_in = testData6[7193];
@(posedge clk);
#1;data_in = testData6[7194];
@(posedge clk);
#1;data_in = testData6[7195];
@(posedge clk);
#1;data_in = testData6[7196];
@(posedge clk);
#1;data_in = testData6[7197];
@(posedge clk);
#1;data_in = testData6[7198];
@(posedge clk);
#1;data_in = testData6[7199];
@(posedge clk);
#1;data_in = testData6[7200];
@(posedge clk);
#1;data_in = testData6[7201];
@(posedge clk);
#1;data_in = testData6[7202];
@(posedge clk);
#1;data_in = testData6[7203];
@(posedge clk);
#1;data_in = testData6[7204];
@(posedge clk);
#1;data_in = testData6[7205];
@(posedge clk);
#1;data_in = testData6[7206];
@(posedge clk);
#1;data_in = testData6[7207];
@(posedge clk);
#1;data_in = testData6[7208];
@(posedge clk);
#1;data_in = testData6[7209];
@(posedge clk);
#1;data_in = testData6[7210];
@(posedge clk);
#1;data_in = testData6[7211];
@(posedge clk);
#1;data_in = testData6[7212];
@(posedge clk);
#1;data_in = testData6[7213];
@(posedge clk);
#1;data_in = testData6[7214];
@(posedge clk);
#1;data_in = testData6[7215];
@(posedge clk);
#1;data_in = testData6[7216];
@(posedge clk);
#1;data_in = testData6[7217];
@(posedge clk);
#1;data_in = testData6[7218];
@(posedge clk);
#1;data_in = testData6[7219];
@(posedge clk);
#1;data_in = testData6[7220];
@(posedge clk);
#1;data_in = testData6[7221];
@(posedge clk);
#1;data_in = testData6[7222];
@(posedge clk);
#1;data_in = testData6[7223];
@(posedge clk);
#1;data_in = testData6[7224];
@(posedge clk);
#1;data_in = testData6[7225];
@(posedge clk);
#1;data_in = testData6[7226];
@(posedge clk);
#1;data_in = testData6[7227];
@(posedge clk);
#1;data_in = testData6[7228];
@(posedge clk);
#1;data_in = testData6[7229];
@(posedge clk);
#1;data_in = testData6[7230];
@(posedge clk);
#1;data_in = testData6[7231];
@(posedge clk);
#1;data_in = testData6[7232];
@(posedge clk);
#1;data_in = testData6[7233];
@(posedge clk);
#1;data_in = testData6[7234];
@(posedge clk);
#1;data_in = testData6[7235];
@(posedge clk);
#1;data_in = testData6[7236];
@(posedge clk);
#1;data_in = testData6[7237];
@(posedge clk);
#1;data_in = testData6[7238];
@(posedge clk);
#1;data_in = testData6[7239];
@(posedge clk);
#1;data_in = testData6[7240];
@(posedge clk);
#1;data_in = testData6[7241];
@(posedge clk);
#1;data_in = testData6[7242];
@(posedge clk);
#1;data_in = testData6[7243];
@(posedge clk);
#1;data_in = testData6[7244];
@(posedge clk);
#1;data_in = testData6[7245];
@(posedge clk);
#1;data_in = testData6[7246];
@(posedge clk);
#1;data_in = testData6[7247];
@(posedge clk);
#1;data_in = testData6[7248];
@(posedge clk);
#1;data_in = testData6[7249];
@(posedge clk);
#1;data_in = testData6[7250];
@(posedge clk);
#1;data_in = testData6[7251];
@(posedge clk);
#1;data_in = testData6[7252];
@(posedge clk);
#1;data_in = testData6[7253];
@(posedge clk);
#1;data_in = testData6[7254];
@(posedge clk);
#1;data_in = testData6[7255];
@(posedge clk);
#1;data_in = testData6[7256];
@(posedge clk);
#1;data_in = testData6[7257];
@(posedge clk);
#1;data_in = testData6[7258];
@(posedge clk);
#1;data_in = testData6[7259];
@(posedge clk);
#1;data_in = testData6[7260];
@(posedge clk);
#1;data_in = testData6[7261];
@(posedge clk);
#1;data_in = testData6[7262];
@(posedge clk);
#1;data_in = testData6[7263];
@(posedge clk);
#1;data_in = testData6[7264];
@(posedge clk);
#1;data_in = testData6[7265];
@(posedge clk);
#1;data_in = testData6[7266];
@(posedge clk);
#1;data_in = testData6[7267];
@(posedge clk);
#1;data_in = testData6[7268];
@(posedge clk);
#1;data_in = testData6[7269];
@(posedge clk);
#1;data_in = testData6[7270];
@(posedge clk);
#1;data_in = testData6[7271];
@(posedge clk);
#1;data_in = testData6[7272];
@(posedge clk);
#1;data_in = testData6[7273];
@(posedge clk);
#1;data_in = testData6[7274];
@(posedge clk);
#1;data_in = testData6[7275];
@(posedge clk);
#1;data_in = testData6[7276];
@(posedge clk);
#1;data_in = testData6[7277];
@(posedge clk);
#1;data_in = testData6[7278];
@(posedge clk);
#1;data_in = testData6[7279];
@(posedge clk);
#1;data_in = testData6[7280];
@(posedge clk);
#1;data_in = testData6[7281];
@(posedge clk);
#1;data_in = testData6[7282];
@(posedge clk);
#1;data_in = testData6[7283];
@(posedge clk);
#1;data_in = testData6[7284];
@(posedge clk);
#1;data_in = testData6[7285];
@(posedge clk);
#1;data_in = testData6[7286];
@(posedge clk);
#1;data_in = testData6[7287];
@(posedge clk);
#1;data_in = testData6[7288];
@(posedge clk);
#1;data_in = testData6[7289];
@(posedge clk);
#1;data_in = testData6[7290];
@(posedge clk);
#1;data_in = testData6[7291];
@(posedge clk);
#1;data_in = testData6[7292];
@(posedge clk);
#1;data_in = testData6[7293];
@(posedge clk);
#1;data_in = testData6[7294];
@(posedge clk);
#1;data_in = testData6[7295];
@(posedge clk);
#1;data_in = testData6[7296];
@(posedge clk);
#1;data_in = testData6[7297];
@(posedge clk);
#1;data_in = testData6[7298];
@(posedge clk);
#1;data_in = testData6[7299];
@(posedge clk);
#1;data_in = testData6[7300];
@(posedge clk);
#1;data_in = testData6[7301];
@(posedge clk);
#1;data_in = testData6[7302];
@(posedge clk);
#1;data_in = testData6[7303];
@(posedge clk);
#1;data_in = testData6[7304];
@(posedge clk);
#1;data_in = testData6[7305];
@(posedge clk);
#1;data_in = testData6[7306];
@(posedge clk);
#1;data_in = testData6[7307];
@(posedge clk);
#1;data_in = testData6[7308];
@(posedge clk);
#1;data_in = testData6[7309];
@(posedge clk);
#1;data_in = testData6[7310];
@(posedge clk);
#1;data_in = testData6[7311];
@(posedge clk);
#1;data_in = testData6[7312];
@(posedge clk);
#1;data_in = testData6[7313];
@(posedge clk);
#1;data_in = testData6[7314];
@(posedge clk);
#1;data_in = testData6[7315];
@(posedge clk);
#1;data_in = testData6[7316];
@(posedge clk);
#1;data_in = testData6[7317];
@(posedge clk);
#1;data_in = testData6[7318];
@(posedge clk);
#1;data_in = testData6[7319];
@(posedge clk);
#1;data_in = testData6[7320];
@(posedge clk);
#1;data_in = testData6[7321];
@(posedge clk);
#1;data_in = testData6[7322];
@(posedge clk);
#1;data_in = testData6[7323];
@(posedge clk);
#1;data_in = testData6[7324];
@(posedge clk);
#1;data_in = testData6[7325];
@(posedge clk);
#1;data_in = testData6[7326];
@(posedge clk);
#1;data_in = testData6[7327];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[7328]; 
@(posedge clk);
#1;data_in = testData6[7329];
@(posedge clk);
#1;data_in = testData6[7330];
@(posedge clk);
#1;data_in = testData6[7331];
@(posedge clk);
#1;data_in = testData6[7332];
@(posedge clk);
#1;data_in = testData6[7333];
@(posedge clk);
#1;data_in = testData6[7334];
@(posedge clk);
#1;data_in = testData6[7335];
@(posedge clk);
#1;data_in = testData6[7336];
@(posedge clk);
#1;data_in = testData6[7337];
@(posedge clk);
#1;data_in = testData6[7338];
@(posedge clk);
#1;data_in = testData6[7339];
@(posedge clk);
#1;data_in = testData6[7340];
@(posedge clk);
#1;data_in = testData6[7341];
@(posedge clk);
#1;data_in = testData6[7342];
@(posedge clk);
#1;data_in = testData6[7343];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[7344];
@(posedge clk);
#1;data_in = testData6[7345];
@(posedge clk);
#1;data_in = testData6[7346];
@(posedge clk);
#1;data_in = testData6[7347];
@(posedge clk);
#1;data_in = testData6[7348];
@(posedge clk);
#1;data_in = testData6[7349];
@(posedge clk);
#1;data_in = testData6[7350];
@(posedge clk);
#1;data_in = testData6[7351];
@(posedge clk);
#1;data_in = testData6[7352];
@(posedge clk);
#1;data_in = testData6[7353];
@(posedge clk);
#1;data_in = testData6[7354];
@(posedge clk);
#1;data_in = testData6[7355];
@(posedge clk);
#1;data_in = testData6[7356];
@(posedge clk);
#1;data_in = testData6[7357];
@(posedge clk);
#1;data_in = testData6[7358];
@(posedge clk);
#1;data_in = testData6[7359];
@(posedge clk);
#1;data_in = testData6[7360];
@(posedge clk);
#1;data_in = testData6[7361];
@(posedge clk);
#1;data_in = testData6[7362];
@(posedge clk);
#1;data_in = testData6[7363];
@(posedge clk);
#1;data_in = testData6[7364];
@(posedge clk);
#1;data_in = testData6[7365];
@(posedge clk);
#1;data_in = testData6[7366];
@(posedge clk);
#1;data_in = testData6[7367];
@(posedge clk);
#1;data_in = testData6[7368];
@(posedge clk);
#1;data_in = testData6[7369];
@(posedge clk);
#1;data_in = testData6[7370];
@(posedge clk);
#1;data_in = testData6[7371];
@(posedge clk);
#1;data_in = testData6[7372];
@(posedge clk);
#1;data_in = testData6[7373];
@(posedge clk);
#1;data_in = testData6[7374];
@(posedge clk);
#1;data_in = testData6[7375];
@(posedge clk);
#1;data_in = testData6[7376];
@(posedge clk);
#1;data_in = testData6[7377];
@(posedge clk);
#1;data_in = testData6[7378];
@(posedge clk);
#1;data_in = testData6[7379];
@(posedge clk);
#1;data_in = testData6[7380];
@(posedge clk);
#1;data_in = testData6[7381];
@(posedge clk);
#1;data_in = testData6[7382];
@(posedge clk);
#1;data_in = testData6[7383];
@(posedge clk);
#1;data_in = testData6[7384];
@(posedge clk);
#1;data_in = testData6[7385];
@(posedge clk);
#1;data_in = testData6[7386];
@(posedge clk);
#1;data_in = testData6[7387];
@(posedge clk);
#1;data_in = testData6[7388];
@(posedge clk);
#1;data_in = testData6[7389];
@(posedge clk);
#1;data_in = testData6[7390];
@(posedge clk);
#1;data_in = testData6[7391];
@(posedge clk);
#1;data_in = testData6[7392];
@(posedge clk);
#1;data_in = testData6[7393];
@(posedge clk);
#1;data_in = testData6[7394];
@(posedge clk);
#1;data_in = testData6[7395];
@(posedge clk);
#1;data_in = testData6[7396];
@(posedge clk);
#1;data_in = testData6[7397];
@(posedge clk);
#1;data_in = testData6[7398];
@(posedge clk);
#1;data_in = testData6[7399];
@(posedge clk);
#1;data_in = testData6[7400];
@(posedge clk);
#1;data_in = testData6[7401];
@(posedge clk);
#1;data_in = testData6[7402];
@(posedge clk);
#1;data_in = testData6[7403];
@(posedge clk);
#1;data_in = testData6[7404];
@(posedge clk);
#1;data_in = testData6[7405];
@(posedge clk);
#1;data_in = testData6[7406];
@(posedge clk);
#1;data_in = testData6[7407];
@(posedge clk);
#1;data_in = testData6[7408];
@(posedge clk);
#1;data_in = testData6[7409];
@(posedge clk);
#1;data_in = testData6[7410];
@(posedge clk);
#1;data_in = testData6[7411];
@(posedge clk);
#1;data_in = testData6[7412];
@(posedge clk);
#1;data_in = testData6[7413];
@(posedge clk);
#1;data_in = testData6[7414];
@(posedge clk);
#1;data_in = testData6[7415];
@(posedge clk);
#1;data_in = testData6[7416];
@(posedge clk);
#1;data_in = testData6[7417];
@(posedge clk);
#1;data_in = testData6[7418];
@(posedge clk);
#1;data_in = testData6[7419];
@(posedge clk);
#1;data_in = testData6[7420];
@(posedge clk);
#1;data_in = testData6[7421];
@(posedge clk);
#1;data_in = testData6[7422];
@(posedge clk);
#1;data_in = testData6[7423];
@(posedge clk);
#1;data_in = testData6[7424];
@(posedge clk);
#1;data_in = testData6[7425];
@(posedge clk);
#1;data_in = testData6[7426];
@(posedge clk);
#1;data_in = testData6[7427];
@(posedge clk);
#1;data_in = testData6[7428];
@(posedge clk);
#1;data_in = testData6[7429];
@(posedge clk);
#1;data_in = testData6[7430];
@(posedge clk);
#1;data_in = testData6[7431];
@(posedge clk);
#1;data_in = testData6[7432];
@(posedge clk);
#1;data_in = testData6[7433];
@(posedge clk);
#1;data_in = testData6[7434];
@(posedge clk);
#1;data_in = testData6[7435];
@(posedge clk);
#1;data_in = testData6[7436];
@(posedge clk);
#1;data_in = testData6[7437];
@(posedge clk);
#1;data_in = testData6[7438];
@(posedge clk);
#1;data_in = testData6[7439];
@(posedge clk);
#1;data_in = testData6[7440];
@(posedge clk);
#1;data_in = testData6[7441];
@(posedge clk);
#1;data_in = testData6[7442];
@(posedge clk);
#1;data_in = testData6[7443];
@(posedge clk);
#1;data_in = testData6[7444];
@(posedge clk);
#1;data_in = testData6[7445];
@(posedge clk);
#1;data_in = testData6[7446];
@(posedge clk);
#1;data_in = testData6[7447];
@(posedge clk);
#1;data_in = testData6[7448];
@(posedge clk);
#1;data_in = testData6[7449];
@(posedge clk);
#1;data_in = testData6[7450];
@(posedge clk);
#1;data_in = testData6[7451];
@(posedge clk);
#1;data_in = testData6[7452];
@(posedge clk);
#1;data_in = testData6[7453];
@(posedge clk);
#1;data_in = testData6[7454];
@(posedge clk);
#1;data_in = testData6[7455];
@(posedge clk);
#1;data_in = testData6[7456];
@(posedge clk);
#1;data_in = testData6[7457];
@(posedge clk);
#1;data_in = testData6[7458];
@(posedge clk);
#1;data_in = testData6[7459];
@(posedge clk);
#1;data_in = testData6[7460];
@(posedge clk);
#1;data_in = testData6[7461];
@(posedge clk);
#1;data_in = testData6[7462];
@(posedge clk);
#1;data_in = testData6[7463];
@(posedge clk);
#1;data_in = testData6[7464];
@(posedge clk);
#1;data_in = testData6[7465];
@(posedge clk);
#1;data_in = testData6[7466];
@(posedge clk);
#1;data_in = testData6[7467];
@(posedge clk);
#1;data_in = testData6[7468];
@(posedge clk);
#1;data_in = testData6[7469];
@(posedge clk);
#1;data_in = testData6[7470];
@(posedge clk);
#1;data_in = testData6[7471];
@(posedge clk);
#1;data_in = testData6[7472];
@(posedge clk);
#1;data_in = testData6[7473];
@(posedge clk);
#1;data_in = testData6[7474];
@(posedge clk);
#1;data_in = testData6[7475];
@(posedge clk);
#1;data_in = testData6[7476];
@(posedge clk);
#1;data_in = testData6[7477];
@(posedge clk);
#1;data_in = testData6[7478];
@(posedge clk);
#1;data_in = testData6[7479];
@(posedge clk);
#1;data_in = testData6[7480];
@(posedge clk);
#1;data_in = testData6[7481];
@(posedge clk);
#1;data_in = testData6[7482];
@(posedge clk);
#1;data_in = testData6[7483];
@(posedge clk);
#1;data_in = testData6[7484];
@(posedge clk);
#1;data_in = testData6[7485];
@(posedge clk);
#1;data_in = testData6[7486];
@(posedge clk);
#1;data_in = testData6[7487];
@(posedge clk);
#1;data_in = testData6[7488];
@(posedge clk);
#1;data_in = testData6[7489];
@(posedge clk);
#1;data_in = testData6[7490];
@(posedge clk);
#1;data_in = testData6[7491];
@(posedge clk);
#1;data_in = testData6[7492];
@(posedge clk);
#1;data_in = testData6[7493];
@(posedge clk);
#1;data_in = testData6[7494];
@(posedge clk);
#1;data_in = testData6[7495];
@(posedge clk);
#1;data_in = testData6[7496];
@(posedge clk);
#1;data_in = testData6[7497];
@(posedge clk);
#1;data_in = testData6[7498];
@(posedge clk);
#1;data_in = testData6[7499];
@(posedge clk);
#1;data_in = testData6[7500];
@(posedge clk);
#1;data_in = testData6[7501];
@(posedge clk);
#1;data_in = testData6[7502];
@(posedge clk);
#1;data_in = testData6[7503];
@(posedge clk);
#1;data_in = testData6[7504];
@(posedge clk);
#1;data_in = testData6[7505];
@(posedge clk);
#1;data_in = testData6[7506];
@(posedge clk);
#1;data_in = testData6[7507];
@(posedge clk);
#1;data_in = testData6[7508];
@(posedge clk);
#1;data_in = testData6[7509];
@(posedge clk);
#1;data_in = testData6[7510];
@(posedge clk);
#1;data_in = testData6[7511];
@(posedge clk);
#1;data_in = testData6[7512];
@(posedge clk);
#1;data_in = testData6[7513];
@(posedge clk);
#1;data_in = testData6[7514];
@(posedge clk);
#1;data_in = testData6[7515];
@(posedge clk);
#1;data_in = testData6[7516];
@(posedge clk);
#1;data_in = testData6[7517];
@(posedge clk);
#1;data_in = testData6[7518];
@(posedge clk);
#1;data_in = testData6[7519];
@(posedge clk);
#1;data_in = testData6[7520];
@(posedge clk);
#1;data_in = testData6[7521];
@(posedge clk);
#1;data_in = testData6[7522];
@(posedge clk);
#1;data_in = testData6[7523];
@(posedge clk);
#1;data_in = testData6[7524];
@(posedge clk);
#1;data_in = testData6[7525];
@(posedge clk);
#1;data_in = testData6[7526];
@(posedge clk);
#1;data_in = testData6[7527];
@(posedge clk);
#1;data_in = testData6[7528];
@(posedge clk);
#1;data_in = testData6[7529];
@(posedge clk);
#1;data_in = testData6[7530];
@(posedge clk);
#1;data_in = testData6[7531];
@(posedge clk);
#1;data_in = testData6[7532];
@(posedge clk);
#1;data_in = testData6[7533];
@(posedge clk);
#1;data_in = testData6[7534];
@(posedge clk);
#1;data_in = testData6[7535];
@(posedge clk);
#1;data_in = testData6[7536];
@(posedge clk);
#1;data_in = testData6[7537];
@(posedge clk);
#1;data_in = testData6[7538];
@(posedge clk);
#1;data_in = testData6[7539];
@(posedge clk);
#1;data_in = testData6[7540];
@(posedge clk);
#1;data_in = testData6[7541];
@(posedge clk);
#1;data_in = testData6[7542];
@(posedge clk);
#1;data_in = testData6[7543];
@(posedge clk);
#1;data_in = testData6[7544];
@(posedge clk);
#1;data_in = testData6[7545];
@(posedge clk);
#1;data_in = testData6[7546];
@(posedge clk);
#1;data_in = testData6[7547];
@(posedge clk);
#1;data_in = testData6[7548];
@(posedge clk);
#1;data_in = testData6[7549];
@(posedge clk);
#1;data_in = testData6[7550];
@(posedge clk);
#1;data_in = testData6[7551];
@(posedge clk);
#1;data_in = testData6[7552];
@(posedge clk);
#1;data_in = testData6[7553];
@(posedge clk);
#1;data_in = testData6[7554];
@(posedge clk);
#1;data_in = testData6[7555];
@(posedge clk);
#1;data_in = testData6[7556];
@(posedge clk);
#1;data_in = testData6[7557];
@(posedge clk);
#1;data_in = testData6[7558];
@(posedge clk);
#1;data_in = testData6[7559];
@(posedge clk);
#1;data_in = testData6[7560];
@(posedge clk);
#1;data_in = testData6[7561];
@(posedge clk);
#1;data_in = testData6[7562];
@(posedge clk);
#1;data_in = testData6[7563];
@(posedge clk);
#1;data_in = testData6[7564];
@(posedge clk);
#1;data_in = testData6[7565];
@(posedge clk);
#1;data_in = testData6[7566];
@(posedge clk);
#1;data_in = testData6[7567];
@(posedge clk);
#1;data_in = testData6[7568];
@(posedge clk);
#1;data_in = testData6[7569];
@(posedge clk);
#1;data_in = testData6[7570];
@(posedge clk);
#1;data_in = testData6[7571];
@(posedge clk);
#1;data_in = testData6[7572];
@(posedge clk);
#1;data_in = testData6[7573];
@(posedge clk);
#1;data_in = testData6[7574];
@(posedge clk);
#1;data_in = testData6[7575];
@(posedge clk);
#1;data_in = testData6[7576];
@(posedge clk);
#1;data_in = testData6[7577];
@(posedge clk);
#1;data_in = testData6[7578];
@(posedge clk);
#1;data_in = testData6[7579];
@(posedge clk);
#1;data_in = testData6[7580];
@(posedge clk);
#1;data_in = testData6[7581];
@(posedge clk);
#1;data_in = testData6[7582];
@(posedge clk);
#1;data_in = testData6[7583];
@(posedge clk);
#1;data_in = testData6[7584];
@(posedge clk);
#1;data_in = testData6[7585];
@(posedge clk);
#1;data_in = testData6[7586];
@(posedge clk);
#1;data_in = testData6[7587];
@(posedge clk);
#1;data_in = testData6[7588];
@(posedge clk);
#1;data_in = testData6[7589];
@(posedge clk);
#1;data_in = testData6[7590];
@(posedge clk);
#1;data_in = testData6[7591];
@(posedge clk);
#1;data_in = testData6[7592];
@(posedge clk);
#1;data_in = testData6[7593];
@(posedge clk);
#1;data_in = testData6[7594];
@(posedge clk);
#1;data_in = testData6[7595];
@(posedge clk);
#1;data_in = testData6[7596];
@(posedge clk);
#1;data_in = testData6[7597];
@(posedge clk);
#1;data_in = testData6[7598];
@(posedge clk);
#1;data_in = testData6[7599];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[7600]; 
@(posedge clk);
#1;data_in = testData6[7601];
@(posedge clk);
#1;data_in = testData6[7602];
@(posedge clk);
#1;data_in = testData6[7603];
@(posedge clk);
#1;data_in = testData6[7604];
@(posedge clk);
#1;data_in = testData6[7605];
@(posedge clk);
#1;data_in = testData6[7606];
@(posedge clk);
#1;data_in = testData6[7607];
@(posedge clk);
#1;data_in = testData6[7608];
@(posedge clk);
#1;data_in = testData6[7609];
@(posedge clk);
#1;data_in = testData6[7610];
@(posedge clk);
#1;data_in = testData6[7611];
@(posedge clk);
#1;data_in = testData6[7612];
@(posedge clk);
#1;data_in = testData6[7613];
@(posedge clk);
#1;data_in = testData6[7614];
@(posedge clk);
#1;data_in = testData6[7615];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[7616];
@(posedge clk);
#1;data_in = testData6[7617];
@(posedge clk);
#1;data_in = testData6[7618];
@(posedge clk);
#1;data_in = testData6[7619];
@(posedge clk);
#1;data_in = testData6[7620];
@(posedge clk);
#1;data_in = testData6[7621];
@(posedge clk);
#1;data_in = testData6[7622];
@(posedge clk);
#1;data_in = testData6[7623];
@(posedge clk);
#1;data_in = testData6[7624];
@(posedge clk);
#1;data_in = testData6[7625];
@(posedge clk);
#1;data_in = testData6[7626];
@(posedge clk);
#1;data_in = testData6[7627];
@(posedge clk);
#1;data_in = testData6[7628];
@(posedge clk);
#1;data_in = testData6[7629];
@(posedge clk);
#1;data_in = testData6[7630];
@(posedge clk);
#1;data_in = testData6[7631];
@(posedge clk);
#1;data_in = testData6[7632];
@(posedge clk);
#1;data_in = testData6[7633];
@(posedge clk);
#1;data_in = testData6[7634];
@(posedge clk);
#1;data_in = testData6[7635];
@(posedge clk);
#1;data_in = testData6[7636];
@(posedge clk);
#1;data_in = testData6[7637];
@(posedge clk);
#1;data_in = testData6[7638];
@(posedge clk);
#1;data_in = testData6[7639];
@(posedge clk);
#1;data_in = testData6[7640];
@(posedge clk);
#1;data_in = testData6[7641];
@(posedge clk);
#1;data_in = testData6[7642];
@(posedge clk);
#1;data_in = testData6[7643];
@(posedge clk);
#1;data_in = testData6[7644];
@(posedge clk);
#1;data_in = testData6[7645];
@(posedge clk);
#1;data_in = testData6[7646];
@(posedge clk);
#1;data_in = testData6[7647];
@(posedge clk);
#1;data_in = testData6[7648];
@(posedge clk);
#1;data_in = testData6[7649];
@(posedge clk);
#1;data_in = testData6[7650];
@(posedge clk);
#1;data_in = testData6[7651];
@(posedge clk);
#1;data_in = testData6[7652];
@(posedge clk);
#1;data_in = testData6[7653];
@(posedge clk);
#1;data_in = testData6[7654];
@(posedge clk);
#1;data_in = testData6[7655];
@(posedge clk);
#1;data_in = testData6[7656];
@(posedge clk);
#1;data_in = testData6[7657];
@(posedge clk);
#1;data_in = testData6[7658];
@(posedge clk);
#1;data_in = testData6[7659];
@(posedge clk);
#1;data_in = testData6[7660];
@(posedge clk);
#1;data_in = testData6[7661];
@(posedge clk);
#1;data_in = testData6[7662];
@(posedge clk);
#1;data_in = testData6[7663];
@(posedge clk);
#1;data_in = testData6[7664];
@(posedge clk);
#1;data_in = testData6[7665];
@(posedge clk);
#1;data_in = testData6[7666];
@(posedge clk);
#1;data_in = testData6[7667];
@(posedge clk);
#1;data_in = testData6[7668];
@(posedge clk);
#1;data_in = testData6[7669];
@(posedge clk);
#1;data_in = testData6[7670];
@(posedge clk);
#1;data_in = testData6[7671];
@(posedge clk);
#1;data_in = testData6[7672];
@(posedge clk);
#1;data_in = testData6[7673];
@(posedge clk);
#1;data_in = testData6[7674];
@(posedge clk);
#1;data_in = testData6[7675];
@(posedge clk);
#1;data_in = testData6[7676];
@(posedge clk);
#1;data_in = testData6[7677];
@(posedge clk);
#1;data_in = testData6[7678];
@(posedge clk);
#1;data_in = testData6[7679];
@(posedge clk);
#1;data_in = testData6[7680];
@(posedge clk);
#1;data_in = testData6[7681];
@(posedge clk);
#1;data_in = testData6[7682];
@(posedge clk);
#1;data_in = testData6[7683];
@(posedge clk);
#1;data_in = testData6[7684];
@(posedge clk);
#1;data_in = testData6[7685];
@(posedge clk);
#1;data_in = testData6[7686];
@(posedge clk);
#1;data_in = testData6[7687];
@(posedge clk);
#1;data_in = testData6[7688];
@(posedge clk);
#1;data_in = testData6[7689];
@(posedge clk);
#1;data_in = testData6[7690];
@(posedge clk);
#1;data_in = testData6[7691];
@(posedge clk);
#1;data_in = testData6[7692];
@(posedge clk);
#1;data_in = testData6[7693];
@(posedge clk);
#1;data_in = testData6[7694];
@(posedge clk);
#1;data_in = testData6[7695];
@(posedge clk);
#1;data_in = testData6[7696];
@(posedge clk);
#1;data_in = testData6[7697];
@(posedge clk);
#1;data_in = testData6[7698];
@(posedge clk);
#1;data_in = testData6[7699];
@(posedge clk);
#1;data_in = testData6[7700];
@(posedge clk);
#1;data_in = testData6[7701];
@(posedge clk);
#1;data_in = testData6[7702];
@(posedge clk);
#1;data_in = testData6[7703];
@(posedge clk);
#1;data_in = testData6[7704];
@(posedge clk);
#1;data_in = testData6[7705];
@(posedge clk);
#1;data_in = testData6[7706];
@(posedge clk);
#1;data_in = testData6[7707];
@(posedge clk);
#1;data_in = testData6[7708];
@(posedge clk);
#1;data_in = testData6[7709];
@(posedge clk);
#1;data_in = testData6[7710];
@(posedge clk);
#1;data_in = testData6[7711];
@(posedge clk);
#1;data_in = testData6[7712];
@(posedge clk);
#1;data_in = testData6[7713];
@(posedge clk);
#1;data_in = testData6[7714];
@(posedge clk);
#1;data_in = testData6[7715];
@(posedge clk);
#1;data_in = testData6[7716];
@(posedge clk);
#1;data_in = testData6[7717];
@(posedge clk);
#1;data_in = testData6[7718];
@(posedge clk);
#1;data_in = testData6[7719];
@(posedge clk);
#1;data_in = testData6[7720];
@(posedge clk);
#1;data_in = testData6[7721];
@(posedge clk);
#1;data_in = testData6[7722];
@(posedge clk);
#1;data_in = testData6[7723];
@(posedge clk);
#1;data_in = testData6[7724];
@(posedge clk);
#1;data_in = testData6[7725];
@(posedge clk);
#1;data_in = testData6[7726];
@(posedge clk);
#1;data_in = testData6[7727];
@(posedge clk);
#1;data_in = testData6[7728];
@(posedge clk);
#1;data_in = testData6[7729];
@(posedge clk);
#1;data_in = testData6[7730];
@(posedge clk);
#1;data_in = testData6[7731];
@(posedge clk);
#1;data_in = testData6[7732];
@(posedge clk);
#1;data_in = testData6[7733];
@(posedge clk);
#1;data_in = testData6[7734];
@(posedge clk);
#1;data_in = testData6[7735];
@(posedge clk);
#1;data_in = testData6[7736];
@(posedge clk);
#1;data_in = testData6[7737];
@(posedge clk);
#1;data_in = testData6[7738];
@(posedge clk);
#1;data_in = testData6[7739];
@(posedge clk);
#1;data_in = testData6[7740];
@(posedge clk);
#1;data_in = testData6[7741];
@(posedge clk);
#1;data_in = testData6[7742];
@(posedge clk);
#1;data_in = testData6[7743];
@(posedge clk);
#1;data_in = testData6[7744];
@(posedge clk);
#1;data_in = testData6[7745];
@(posedge clk);
#1;data_in = testData6[7746];
@(posedge clk);
#1;data_in = testData6[7747];
@(posedge clk);
#1;data_in = testData6[7748];
@(posedge clk);
#1;data_in = testData6[7749];
@(posedge clk);
#1;data_in = testData6[7750];
@(posedge clk);
#1;data_in = testData6[7751];
@(posedge clk);
#1;data_in = testData6[7752];
@(posedge clk);
#1;data_in = testData6[7753];
@(posedge clk);
#1;data_in = testData6[7754];
@(posedge clk);
#1;data_in = testData6[7755];
@(posedge clk);
#1;data_in = testData6[7756];
@(posedge clk);
#1;data_in = testData6[7757];
@(posedge clk);
#1;data_in = testData6[7758];
@(posedge clk);
#1;data_in = testData6[7759];
@(posedge clk);
#1;data_in = testData6[7760];
@(posedge clk);
#1;data_in = testData6[7761];
@(posedge clk);
#1;data_in = testData6[7762];
@(posedge clk);
#1;data_in = testData6[7763];
@(posedge clk);
#1;data_in = testData6[7764];
@(posedge clk);
#1;data_in = testData6[7765];
@(posedge clk);
#1;data_in = testData6[7766];
@(posedge clk);
#1;data_in = testData6[7767];
@(posedge clk);
#1;data_in = testData6[7768];
@(posedge clk);
#1;data_in = testData6[7769];
@(posedge clk);
#1;data_in = testData6[7770];
@(posedge clk);
#1;data_in = testData6[7771];
@(posedge clk);
#1;data_in = testData6[7772];
@(posedge clk);
#1;data_in = testData6[7773];
@(posedge clk);
#1;data_in = testData6[7774];
@(posedge clk);
#1;data_in = testData6[7775];
@(posedge clk);
#1;data_in = testData6[7776];
@(posedge clk);
#1;data_in = testData6[7777];
@(posedge clk);
#1;data_in = testData6[7778];
@(posedge clk);
#1;data_in = testData6[7779];
@(posedge clk);
#1;data_in = testData6[7780];
@(posedge clk);
#1;data_in = testData6[7781];
@(posedge clk);
#1;data_in = testData6[7782];
@(posedge clk);
#1;data_in = testData6[7783];
@(posedge clk);
#1;data_in = testData6[7784];
@(posedge clk);
#1;data_in = testData6[7785];
@(posedge clk);
#1;data_in = testData6[7786];
@(posedge clk);
#1;data_in = testData6[7787];
@(posedge clk);
#1;data_in = testData6[7788];
@(posedge clk);
#1;data_in = testData6[7789];
@(posedge clk);
#1;data_in = testData6[7790];
@(posedge clk);
#1;data_in = testData6[7791];
@(posedge clk);
#1;data_in = testData6[7792];
@(posedge clk);
#1;data_in = testData6[7793];
@(posedge clk);
#1;data_in = testData6[7794];
@(posedge clk);
#1;data_in = testData6[7795];
@(posedge clk);
#1;data_in = testData6[7796];
@(posedge clk);
#1;data_in = testData6[7797];
@(posedge clk);
#1;data_in = testData6[7798];
@(posedge clk);
#1;data_in = testData6[7799];
@(posedge clk);
#1;data_in = testData6[7800];
@(posedge clk);
#1;data_in = testData6[7801];
@(posedge clk);
#1;data_in = testData6[7802];
@(posedge clk);
#1;data_in = testData6[7803];
@(posedge clk);
#1;data_in = testData6[7804];
@(posedge clk);
#1;data_in = testData6[7805];
@(posedge clk);
#1;data_in = testData6[7806];
@(posedge clk);
#1;data_in = testData6[7807];
@(posedge clk);
#1;data_in = testData6[7808];
@(posedge clk);
#1;data_in = testData6[7809];
@(posedge clk);
#1;data_in = testData6[7810];
@(posedge clk);
#1;data_in = testData6[7811];
@(posedge clk);
#1;data_in = testData6[7812];
@(posedge clk);
#1;data_in = testData6[7813];
@(posedge clk);
#1;data_in = testData6[7814];
@(posedge clk);
#1;data_in = testData6[7815];
@(posedge clk);
#1;data_in = testData6[7816];
@(posedge clk);
#1;data_in = testData6[7817];
@(posedge clk);
#1;data_in = testData6[7818];
@(posedge clk);
#1;data_in = testData6[7819];
@(posedge clk);
#1;data_in = testData6[7820];
@(posedge clk);
#1;data_in = testData6[7821];
@(posedge clk);
#1;data_in = testData6[7822];
@(posedge clk);
#1;data_in = testData6[7823];
@(posedge clk);
#1;data_in = testData6[7824];
@(posedge clk);
#1;data_in = testData6[7825];
@(posedge clk);
#1;data_in = testData6[7826];
@(posedge clk);
#1;data_in = testData6[7827];
@(posedge clk);
#1;data_in = testData6[7828];
@(posedge clk);
#1;data_in = testData6[7829];
@(posedge clk);
#1;data_in = testData6[7830];
@(posedge clk);
#1;data_in = testData6[7831];
@(posedge clk);
#1;data_in = testData6[7832];
@(posedge clk);
#1;data_in = testData6[7833];
@(posedge clk);
#1;data_in = testData6[7834];
@(posedge clk);
#1;data_in = testData6[7835];
@(posedge clk);
#1;data_in = testData6[7836];
@(posedge clk);
#1;data_in = testData6[7837];
@(posedge clk);
#1;data_in = testData6[7838];
@(posedge clk);
#1;data_in = testData6[7839];
@(posedge clk);
#1;data_in = testData6[7840];
@(posedge clk);
#1;data_in = testData6[7841];
@(posedge clk);
#1;data_in = testData6[7842];
@(posedge clk);
#1;data_in = testData6[7843];
@(posedge clk);
#1;data_in = testData6[7844];
@(posedge clk);
#1;data_in = testData6[7845];
@(posedge clk);
#1;data_in = testData6[7846];
@(posedge clk);
#1;data_in = testData6[7847];
@(posedge clk);
#1;data_in = testData6[7848];
@(posedge clk);
#1;data_in = testData6[7849];
@(posedge clk);
#1;data_in = testData6[7850];
@(posedge clk);
#1;data_in = testData6[7851];
@(posedge clk);
#1;data_in = testData6[7852];
@(posedge clk);
#1;data_in = testData6[7853];
@(posedge clk);
#1;data_in = testData6[7854];
@(posedge clk);
#1;data_in = testData6[7855];
@(posedge clk);
#1;data_in = testData6[7856];
@(posedge clk);
#1;data_in = testData6[7857];
@(posedge clk);
#1;data_in = testData6[7858];
@(posedge clk);
#1;data_in = testData6[7859];
@(posedge clk);
#1;data_in = testData6[7860];
@(posedge clk);
#1;data_in = testData6[7861];
@(posedge clk);
#1;data_in = testData6[7862];
@(posedge clk);
#1;data_in = testData6[7863];
@(posedge clk);
#1;data_in = testData6[7864];
@(posedge clk);
#1;data_in = testData6[7865];
@(posedge clk);
#1;data_in = testData6[7866];
@(posedge clk);
#1;data_in = testData6[7867];
@(posedge clk);
#1;data_in = testData6[7868];
@(posedge clk);
#1;data_in = testData6[7869];
@(posedge clk);
#1;data_in = testData6[7870];
@(posedge clk);
#1;data_in = testData6[7871];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[7872]; 
@(posedge clk);
#1;data_in = testData6[7873];
@(posedge clk);
#1;data_in = testData6[7874];
@(posedge clk);
#1;data_in = testData6[7875];
@(posedge clk);
#1;data_in = testData6[7876];
@(posedge clk);
#1;data_in = testData6[7877];
@(posedge clk);
#1;data_in = testData6[7878];
@(posedge clk);
#1;data_in = testData6[7879];
@(posedge clk);
#1;data_in = testData6[7880];
@(posedge clk);
#1;data_in = testData6[7881];
@(posedge clk);
#1;data_in = testData6[7882];
@(posedge clk);
#1;data_in = testData6[7883];
@(posedge clk);
#1;data_in = testData6[7884];
@(posedge clk);
#1;data_in = testData6[7885];
@(posedge clk);
#1;data_in = testData6[7886];
@(posedge clk);
#1;data_in = testData6[7887];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[7888];
@(posedge clk);
#1;data_in = testData6[7889];
@(posedge clk);
#1;data_in = testData6[7890];
@(posedge clk);
#1;data_in = testData6[7891];
@(posedge clk);
#1;data_in = testData6[7892];
@(posedge clk);
#1;data_in = testData6[7893];
@(posedge clk);
#1;data_in = testData6[7894];
@(posedge clk);
#1;data_in = testData6[7895];
@(posedge clk);
#1;data_in = testData6[7896];
@(posedge clk);
#1;data_in = testData6[7897];
@(posedge clk);
#1;data_in = testData6[7898];
@(posedge clk);
#1;data_in = testData6[7899];
@(posedge clk);
#1;data_in = testData6[7900];
@(posedge clk);
#1;data_in = testData6[7901];
@(posedge clk);
#1;data_in = testData6[7902];
@(posedge clk);
#1;data_in = testData6[7903];
@(posedge clk);
#1;data_in = testData6[7904];
@(posedge clk);
#1;data_in = testData6[7905];
@(posedge clk);
#1;data_in = testData6[7906];
@(posedge clk);
#1;data_in = testData6[7907];
@(posedge clk);
#1;data_in = testData6[7908];
@(posedge clk);
#1;data_in = testData6[7909];
@(posedge clk);
#1;data_in = testData6[7910];
@(posedge clk);
#1;data_in = testData6[7911];
@(posedge clk);
#1;data_in = testData6[7912];
@(posedge clk);
#1;data_in = testData6[7913];
@(posedge clk);
#1;data_in = testData6[7914];
@(posedge clk);
#1;data_in = testData6[7915];
@(posedge clk);
#1;data_in = testData6[7916];
@(posedge clk);
#1;data_in = testData6[7917];
@(posedge clk);
#1;data_in = testData6[7918];
@(posedge clk);
#1;data_in = testData6[7919];
@(posedge clk);
#1;data_in = testData6[7920];
@(posedge clk);
#1;data_in = testData6[7921];
@(posedge clk);
#1;data_in = testData6[7922];
@(posedge clk);
#1;data_in = testData6[7923];
@(posedge clk);
#1;data_in = testData6[7924];
@(posedge clk);
#1;data_in = testData6[7925];
@(posedge clk);
#1;data_in = testData6[7926];
@(posedge clk);
#1;data_in = testData6[7927];
@(posedge clk);
#1;data_in = testData6[7928];
@(posedge clk);
#1;data_in = testData6[7929];
@(posedge clk);
#1;data_in = testData6[7930];
@(posedge clk);
#1;data_in = testData6[7931];
@(posedge clk);
#1;data_in = testData6[7932];
@(posedge clk);
#1;data_in = testData6[7933];
@(posedge clk);
#1;data_in = testData6[7934];
@(posedge clk);
#1;data_in = testData6[7935];
@(posedge clk);
#1;data_in = testData6[7936];
@(posedge clk);
#1;data_in = testData6[7937];
@(posedge clk);
#1;data_in = testData6[7938];
@(posedge clk);
#1;data_in = testData6[7939];
@(posedge clk);
#1;data_in = testData6[7940];
@(posedge clk);
#1;data_in = testData6[7941];
@(posedge clk);
#1;data_in = testData6[7942];
@(posedge clk);
#1;data_in = testData6[7943];
@(posedge clk);
#1;data_in = testData6[7944];
@(posedge clk);
#1;data_in = testData6[7945];
@(posedge clk);
#1;data_in = testData6[7946];
@(posedge clk);
#1;data_in = testData6[7947];
@(posedge clk);
#1;data_in = testData6[7948];
@(posedge clk);
#1;data_in = testData6[7949];
@(posedge clk);
#1;data_in = testData6[7950];
@(posedge clk);
#1;data_in = testData6[7951];
@(posedge clk);
#1;data_in = testData6[7952];
@(posedge clk);
#1;data_in = testData6[7953];
@(posedge clk);
#1;data_in = testData6[7954];
@(posedge clk);
#1;data_in = testData6[7955];
@(posedge clk);
#1;data_in = testData6[7956];
@(posedge clk);
#1;data_in = testData6[7957];
@(posedge clk);
#1;data_in = testData6[7958];
@(posedge clk);
#1;data_in = testData6[7959];
@(posedge clk);
#1;data_in = testData6[7960];
@(posedge clk);
#1;data_in = testData6[7961];
@(posedge clk);
#1;data_in = testData6[7962];
@(posedge clk);
#1;data_in = testData6[7963];
@(posedge clk);
#1;data_in = testData6[7964];
@(posedge clk);
#1;data_in = testData6[7965];
@(posedge clk);
#1;data_in = testData6[7966];
@(posedge clk);
#1;data_in = testData6[7967];
@(posedge clk);
#1;data_in = testData6[7968];
@(posedge clk);
#1;data_in = testData6[7969];
@(posedge clk);
#1;data_in = testData6[7970];
@(posedge clk);
#1;data_in = testData6[7971];
@(posedge clk);
#1;data_in = testData6[7972];
@(posedge clk);
#1;data_in = testData6[7973];
@(posedge clk);
#1;data_in = testData6[7974];
@(posedge clk);
#1;data_in = testData6[7975];
@(posedge clk);
#1;data_in = testData6[7976];
@(posedge clk);
#1;data_in = testData6[7977];
@(posedge clk);
#1;data_in = testData6[7978];
@(posedge clk);
#1;data_in = testData6[7979];
@(posedge clk);
#1;data_in = testData6[7980];
@(posedge clk);
#1;data_in = testData6[7981];
@(posedge clk);
#1;data_in = testData6[7982];
@(posedge clk);
#1;data_in = testData6[7983];
@(posedge clk);
#1;data_in = testData6[7984];
@(posedge clk);
#1;data_in = testData6[7985];
@(posedge clk);
#1;data_in = testData6[7986];
@(posedge clk);
#1;data_in = testData6[7987];
@(posedge clk);
#1;data_in = testData6[7988];
@(posedge clk);
#1;data_in = testData6[7989];
@(posedge clk);
#1;data_in = testData6[7990];
@(posedge clk);
#1;data_in = testData6[7991];
@(posedge clk);
#1;data_in = testData6[7992];
@(posedge clk);
#1;data_in = testData6[7993];
@(posedge clk);
#1;data_in = testData6[7994];
@(posedge clk);
#1;data_in = testData6[7995];
@(posedge clk);
#1;data_in = testData6[7996];
@(posedge clk);
#1;data_in = testData6[7997];
@(posedge clk);
#1;data_in = testData6[7998];
@(posedge clk);
#1;data_in = testData6[7999];
@(posedge clk);
#1;data_in = testData6[8000];
@(posedge clk);
#1;data_in = testData6[8001];
@(posedge clk);
#1;data_in = testData6[8002];
@(posedge clk);
#1;data_in = testData6[8003];
@(posedge clk);
#1;data_in = testData6[8004];
@(posedge clk);
#1;data_in = testData6[8005];
@(posedge clk);
#1;data_in = testData6[8006];
@(posedge clk);
#1;data_in = testData6[8007];
@(posedge clk);
#1;data_in = testData6[8008];
@(posedge clk);
#1;data_in = testData6[8009];
@(posedge clk);
#1;data_in = testData6[8010];
@(posedge clk);
#1;data_in = testData6[8011];
@(posedge clk);
#1;data_in = testData6[8012];
@(posedge clk);
#1;data_in = testData6[8013];
@(posedge clk);
#1;data_in = testData6[8014];
@(posedge clk);
#1;data_in = testData6[8015];
@(posedge clk);
#1;data_in = testData6[8016];
@(posedge clk);
#1;data_in = testData6[8017];
@(posedge clk);
#1;data_in = testData6[8018];
@(posedge clk);
#1;data_in = testData6[8019];
@(posedge clk);
#1;data_in = testData6[8020];
@(posedge clk);
#1;data_in = testData6[8021];
@(posedge clk);
#1;data_in = testData6[8022];
@(posedge clk);
#1;data_in = testData6[8023];
@(posedge clk);
#1;data_in = testData6[8024];
@(posedge clk);
#1;data_in = testData6[8025];
@(posedge clk);
#1;data_in = testData6[8026];
@(posedge clk);
#1;data_in = testData6[8027];
@(posedge clk);
#1;data_in = testData6[8028];
@(posedge clk);
#1;data_in = testData6[8029];
@(posedge clk);
#1;data_in = testData6[8030];
@(posedge clk);
#1;data_in = testData6[8031];
@(posedge clk);
#1;data_in = testData6[8032];
@(posedge clk);
#1;data_in = testData6[8033];
@(posedge clk);
#1;data_in = testData6[8034];
@(posedge clk);
#1;data_in = testData6[8035];
@(posedge clk);
#1;data_in = testData6[8036];
@(posedge clk);
#1;data_in = testData6[8037];
@(posedge clk);
#1;data_in = testData6[8038];
@(posedge clk);
#1;data_in = testData6[8039];
@(posedge clk);
#1;data_in = testData6[8040];
@(posedge clk);
#1;data_in = testData6[8041];
@(posedge clk);
#1;data_in = testData6[8042];
@(posedge clk);
#1;data_in = testData6[8043];
@(posedge clk);
#1;data_in = testData6[8044];
@(posedge clk);
#1;data_in = testData6[8045];
@(posedge clk);
#1;data_in = testData6[8046];
@(posedge clk);
#1;data_in = testData6[8047];
@(posedge clk);
#1;data_in = testData6[8048];
@(posedge clk);
#1;data_in = testData6[8049];
@(posedge clk);
#1;data_in = testData6[8050];
@(posedge clk);
#1;data_in = testData6[8051];
@(posedge clk);
#1;data_in = testData6[8052];
@(posedge clk);
#1;data_in = testData6[8053];
@(posedge clk);
#1;data_in = testData6[8054];
@(posedge clk);
#1;data_in = testData6[8055];
@(posedge clk);
#1;data_in = testData6[8056];
@(posedge clk);
#1;data_in = testData6[8057];
@(posedge clk);
#1;data_in = testData6[8058];
@(posedge clk);
#1;data_in = testData6[8059];
@(posedge clk);
#1;data_in = testData6[8060];
@(posedge clk);
#1;data_in = testData6[8061];
@(posedge clk);
#1;data_in = testData6[8062];
@(posedge clk);
#1;data_in = testData6[8063];
@(posedge clk);
#1;data_in = testData6[8064];
@(posedge clk);
#1;data_in = testData6[8065];
@(posedge clk);
#1;data_in = testData6[8066];
@(posedge clk);
#1;data_in = testData6[8067];
@(posedge clk);
#1;data_in = testData6[8068];
@(posedge clk);
#1;data_in = testData6[8069];
@(posedge clk);
#1;data_in = testData6[8070];
@(posedge clk);
#1;data_in = testData6[8071];
@(posedge clk);
#1;data_in = testData6[8072];
@(posedge clk);
#1;data_in = testData6[8073];
@(posedge clk);
#1;data_in = testData6[8074];
@(posedge clk);
#1;data_in = testData6[8075];
@(posedge clk);
#1;data_in = testData6[8076];
@(posedge clk);
#1;data_in = testData6[8077];
@(posedge clk);
#1;data_in = testData6[8078];
@(posedge clk);
#1;data_in = testData6[8079];
@(posedge clk);
#1;data_in = testData6[8080];
@(posedge clk);
#1;data_in = testData6[8081];
@(posedge clk);
#1;data_in = testData6[8082];
@(posedge clk);
#1;data_in = testData6[8083];
@(posedge clk);
#1;data_in = testData6[8084];
@(posedge clk);
#1;data_in = testData6[8085];
@(posedge clk);
#1;data_in = testData6[8086];
@(posedge clk);
#1;data_in = testData6[8087];
@(posedge clk);
#1;data_in = testData6[8088];
@(posedge clk);
#1;data_in = testData6[8089];
@(posedge clk);
#1;data_in = testData6[8090];
@(posedge clk);
#1;data_in = testData6[8091];
@(posedge clk);
#1;data_in = testData6[8092];
@(posedge clk);
#1;data_in = testData6[8093];
@(posedge clk);
#1;data_in = testData6[8094];
@(posedge clk);
#1;data_in = testData6[8095];
@(posedge clk);
#1;data_in = testData6[8096];
@(posedge clk);
#1;data_in = testData6[8097];
@(posedge clk);
#1;data_in = testData6[8098];
@(posedge clk);
#1;data_in = testData6[8099];
@(posedge clk);
#1;data_in = testData6[8100];
@(posedge clk);
#1;data_in = testData6[8101];
@(posedge clk);
#1;data_in = testData6[8102];
@(posedge clk);
#1;data_in = testData6[8103];
@(posedge clk);
#1;data_in = testData6[8104];
@(posedge clk);
#1;data_in = testData6[8105];
@(posedge clk);
#1;data_in = testData6[8106];
@(posedge clk);
#1;data_in = testData6[8107];
@(posedge clk);
#1;data_in = testData6[8108];
@(posedge clk);
#1;data_in = testData6[8109];
@(posedge clk);
#1;data_in = testData6[8110];
@(posedge clk);
#1;data_in = testData6[8111];
@(posedge clk);
#1;data_in = testData6[8112];
@(posedge clk);
#1;data_in = testData6[8113];
@(posedge clk);
#1;data_in = testData6[8114];
@(posedge clk);
#1;data_in = testData6[8115];
@(posedge clk);
#1;data_in = testData6[8116];
@(posedge clk);
#1;data_in = testData6[8117];
@(posedge clk);
#1;data_in = testData6[8118];
@(posedge clk);
#1;data_in = testData6[8119];
@(posedge clk);
#1;data_in = testData6[8120];
@(posedge clk);
#1;data_in = testData6[8121];
@(posedge clk);
#1;data_in = testData6[8122];
@(posedge clk);
#1;data_in = testData6[8123];
@(posedge clk);
#1;data_in = testData6[8124];
@(posedge clk);
#1;data_in = testData6[8125];
@(posedge clk);
#1;data_in = testData6[8126];
@(posedge clk);
#1;data_in = testData6[8127];
@(posedge clk);
#1;data_in = testData6[8128];
@(posedge clk);
#1;data_in = testData6[8129];
@(posedge clk);
#1;data_in = testData6[8130];
@(posedge clk);
#1;data_in = testData6[8131];
@(posedge clk);
#1;data_in = testData6[8132];
@(posedge clk);
#1;data_in = testData6[8133];
@(posedge clk);
#1;data_in = testData6[8134];
@(posedge clk);
#1;data_in = testData6[8135];
@(posedge clk);
#1;data_in = testData6[8136];
@(posedge clk);
#1;data_in = testData6[8137];
@(posedge clk);
#1;data_in = testData6[8138];
@(posedge clk);
#1;data_in = testData6[8139];
@(posedge clk);
#1;data_in = testData6[8140];
@(posedge clk);
#1;data_in = testData6[8141];
@(posedge clk);
#1;data_in = testData6[8142];
@(posedge clk);
#1;data_in = testData6[8143];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[8144]; 
@(posedge clk);
#1;data_in = testData6[8145];
@(posedge clk);
#1;data_in = testData6[8146];
@(posedge clk);
#1;data_in = testData6[8147];
@(posedge clk);
#1;data_in = testData6[8148];
@(posedge clk);
#1;data_in = testData6[8149];
@(posedge clk);
#1;data_in = testData6[8150];
@(posedge clk);
#1;data_in = testData6[8151];
@(posedge clk);
#1;data_in = testData6[8152];
@(posedge clk);
#1;data_in = testData6[8153];
@(posedge clk);
#1;data_in = testData6[8154];
@(posedge clk);
#1;data_in = testData6[8155];
@(posedge clk);
#1;data_in = testData6[8156];
@(posedge clk);
#1;data_in = testData6[8157];
@(posedge clk);
#1;data_in = testData6[8158];
@(posedge clk);
#1;data_in = testData6[8159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[8160];
@(posedge clk);
#1;data_in = testData6[8161];
@(posedge clk);
#1;data_in = testData6[8162];
@(posedge clk);
#1;data_in = testData6[8163];
@(posedge clk);
#1;data_in = testData6[8164];
@(posedge clk);
#1;data_in = testData6[8165];
@(posedge clk);
#1;data_in = testData6[8166];
@(posedge clk);
#1;data_in = testData6[8167];
@(posedge clk);
#1;data_in = testData6[8168];
@(posedge clk);
#1;data_in = testData6[8169];
@(posedge clk);
#1;data_in = testData6[8170];
@(posedge clk);
#1;data_in = testData6[8171];
@(posedge clk);
#1;data_in = testData6[8172];
@(posedge clk);
#1;data_in = testData6[8173];
@(posedge clk);
#1;data_in = testData6[8174];
@(posedge clk);
#1;data_in = testData6[8175];
@(posedge clk);
#1;data_in = testData6[8176];
@(posedge clk);
#1;data_in = testData6[8177];
@(posedge clk);
#1;data_in = testData6[8178];
@(posedge clk);
#1;data_in = testData6[8179];
@(posedge clk);
#1;data_in = testData6[8180];
@(posedge clk);
#1;data_in = testData6[8181];
@(posedge clk);
#1;data_in = testData6[8182];
@(posedge clk);
#1;data_in = testData6[8183];
@(posedge clk);
#1;data_in = testData6[8184];
@(posedge clk);
#1;data_in = testData6[8185];
@(posedge clk);
#1;data_in = testData6[8186];
@(posedge clk);
#1;data_in = testData6[8187];
@(posedge clk);
#1;data_in = testData6[8188];
@(posedge clk);
#1;data_in = testData6[8189];
@(posedge clk);
#1;data_in = testData6[8190];
@(posedge clk);
#1;data_in = testData6[8191];
@(posedge clk);
#1;data_in = testData6[8192];
@(posedge clk);
#1;data_in = testData6[8193];
@(posedge clk);
#1;data_in = testData6[8194];
@(posedge clk);
#1;data_in = testData6[8195];
@(posedge clk);
#1;data_in = testData6[8196];
@(posedge clk);
#1;data_in = testData6[8197];
@(posedge clk);
#1;data_in = testData6[8198];
@(posedge clk);
#1;data_in = testData6[8199];
@(posedge clk);
#1;data_in = testData6[8200];
@(posedge clk);
#1;data_in = testData6[8201];
@(posedge clk);
#1;data_in = testData6[8202];
@(posedge clk);
#1;data_in = testData6[8203];
@(posedge clk);
#1;data_in = testData6[8204];
@(posedge clk);
#1;data_in = testData6[8205];
@(posedge clk);
#1;data_in = testData6[8206];
@(posedge clk);
#1;data_in = testData6[8207];
@(posedge clk);
#1;data_in = testData6[8208];
@(posedge clk);
#1;data_in = testData6[8209];
@(posedge clk);
#1;data_in = testData6[8210];
@(posedge clk);
#1;data_in = testData6[8211];
@(posedge clk);
#1;data_in = testData6[8212];
@(posedge clk);
#1;data_in = testData6[8213];
@(posedge clk);
#1;data_in = testData6[8214];
@(posedge clk);
#1;data_in = testData6[8215];
@(posedge clk);
#1;data_in = testData6[8216];
@(posedge clk);
#1;data_in = testData6[8217];
@(posedge clk);
#1;data_in = testData6[8218];
@(posedge clk);
#1;data_in = testData6[8219];
@(posedge clk);
#1;data_in = testData6[8220];
@(posedge clk);
#1;data_in = testData6[8221];
@(posedge clk);
#1;data_in = testData6[8222];
@(posedge clk);
#1;data_in = testData6[8223];
@(posedge clk);
#1;data_in = testData6[8224];
@(posedge clk);
#1;data_in = testData6[8225];
@(posedge clk);
#1;data_in = testData6[8226];
@(posedge clk);
#1;data_in = testData6[8227];
@(posedge clk);
#1;data_in = testData6[8228];
@(posedge clk);
#1;data_in = testData6[8229];
@(posedge clk);
#1;data_in = testData6[8230];
@(posedge clk);
#1;data_in = testData6[8231];
@(posedge clk);
#1;data_in = testData6[8232];
@(posedge clk);
#1;data_in = testData6[8233];
@(posedge clk);
#1;data_in = testData6[8234];
@(posedge clk);
#1;data_in = testData6[8235];
@(posedge clk);
#1;data_in = testData6[8236];
@(posedge clk);
#1;data_in = testData6[8237];
@(posedge clk);
#1;data_in = testData6[8238];
@(posedge clk);
#1;data_in = testData6[8239];
@(posedge clk);
#1;data_in = testData6[8240];
@(posedge clk);
#1;data_in = testData6[8241];
@(posedge clk);
#1;data_in = testData6[8242];
@(posedge clk);
#1;data_in = testData6[8243];
@(posedge clk);
#1;data_in = testData6[8244];
@(posedge clk);
#1;data_in = testData6[8245];
@(posedge clk);
#1;data_in = testData6[8246];
@(posedge clk);
#1;data_in = testData6[8247];
@(posedge clk);
#1;data_in = testData6[8248];
@(posedge clk);
#1;data_in = testData6[8249];
@(posedge clk);
#1;data_in = testData6[8250];
@(posedge clk);
#1;data_in = testData6[8251];
@(posedge clk);
#1;data_in = testData6[8252];
@(posedge clk);
#1;data_in = testData6[8253];
@(posedge clk);
#1;data_in = testData6[8254];
@(posedge clk);
#1;data_in = testData6[8255];
@(posedge clk);
#1;data_in = testData6[8256];
@(posedge clk);
#1;data_in = testData6[8257];
@(posedge clk);
#1;data_in = testData6[8258];
@(posedge clk);
#1;data_in = testData6[8259];
@(posedge clk);
#1;data_in = testData6[8260];
@(posedge clk);
#1;data_in = testData6[8261];
@(posedge clk);
#1;data_in = testData6[8262];
@(posedge clk);
#1;data_in = testData6[8263];
@(posedge clk);
#1;data_in = testData6[8264];
@(posedge clk);
#1;data_in = testData6[8265];
@(posedge clk);
#1;data_in = testData6[8266];
@(posedge clk);
#1;data_in = testData6[8267];
@(posedge clk);
#1;data_in = testData6[8268];
@(posedge clk);
#1;data_in = testData6[8269];
@(posedge clk);
#1;data_in = testData6[8270];
@(posedge clk);
#1;data_in = testData6[8271];
@(posedge clk);
#1;data_in = testData6[8272];
@(posedge clk);
#1;data_in = testData6[8273];
@(posedge clk);
#1;data_in = testData6[8274];
@(posedge clk);
#1;data_in = testData6[8275];
@(posedge clk);
#1;data_in = testData6[8276];
@(posedge clk);
#1;data_in = testData6[8277];
@(posedge clk);
#1;data_in = testData6[8278];
@(posedge clk);
#1;data_in = testData6[8279];
@(posedge clk);
#1;data_in = testData6[8280];
@(posedge clk);
#1;data_in = testData6[8281];
@(posedge clk);
#1;data_in = testData6[8282];
@(posedge clk);
#1;data_in = testData6[8283];
@(posedge clk);
#1;data_in = testData6[8284];
@(posedge clk);
#1;data_in = testData6[8285];
@(posedge clk);
#1;data_in = testData6[8286];
@(posedge clk);
#1;data_in = testData6[8287];
@(posedge clk);
#1;data_in = testData6[8288];
@(posedge clk);
#1;data_in = testData6[8289];
@(posedge clk);
#1;data_in = testData6[8290];
@(posedge clk);
#1;data_in = testData6[8291];
@(posedge clk);
#1;data_in = testData6[8292];
@(posedge clk);
#1;data_in = testData6[8293];
@(posedge clk);
#1;data_in = testData6[8294];
@(posedge clk);
#1;data_in = testData6[8295];
@(posedge clk);
#1;data_in = testData6[8296];
@(posedge clk);
#1;data_in = testData6[8297];
@(posedge clk);
#1;data_in = testData6[8298];
@(posedge clk);
#1;data_in = testData6[8299];
@(posedge clk);
#1;data_in = testData6[8300];
@(posedge clk);
#1;data_in = testData6[8301];
@(posedge clk);
#1;data_in = testData6[8302];
@(posedge clk);
#1;data_in = testData6[8303];
@(posedge clk);
#1;data_in = testData6[8304];
@(posedge clk);
#1;data_in = testData6[8305];
@(posedge clk);
#1;data_in = testData6[8306];
@(posedge clk);
#1;data_in = testData6[8307];
@(posedge clk);
#1;data_in = testData6[8308];
@(posedge clk);
#1;data_in = testData6[8309];
@(posedge clk);
#1;data_in = testData6[8310];
@(posedge clk);
#1;data_in = testData6[8311];
@(posedge clk);
#1;data_in = testData6[8312];
@(posedge clk);
#1;data_in = testData6[8313];
@(posedge clk);
#1;data_in = testData6[8314];
@(posedge clk);
#1;data_in = testData6[8315];
@(posedge clk);
#1;data_in = testData6[8316];
@(posedge clk);
#1;data_in = testData6[8317];
@(posedge clk);
#1;data_in = testData6[8318];
@(posedge clk);
#1;data_in = testData6[8319];
@(posedge clk);
#1;data_in = testData6[8320];
@(posedge clk);
#1;data_in = testData6[8321];
@(posedge clk);
#1;data_in = testData6[8322];
@(posedge clk);
#1;data_in = testData6[8323];
@(posedge clk);
#1;data_in = testData6[8324];
@(posedge clk);
#1;data_in = testData6[8325];
@(posedge clk);
#1;data_in = testData6[8326];
@(posedge clk);
#1;data_in = testData6[8327];
@(posedge clk);
#1;data_in = testData6[8328];
@(posedge clk);
#1;data_in = testData6[8329];
@(posedge clk);
#1;data_in = testData6[8330];
@(posedge clk);
#1;data_in = testData6[8331];
@(posedge clk);
#1;data_in = testData6[8332];
@(posedge clk);
#1;data_in = testData6[8333];
@(posedge clk);
#1;data_in = testData6[8334];
@(posedge clk);
#1;data_in = testData6[8335];
@(posedge clk);
#1;data_in = testData6[8336];
@(posedge clk);
#1;data_in = testData6[8337];
@(posedge clk);
#1;data_in = testData6[8338];
@(posedge clk);
#1;data_in = testData6[8339];
@(posedge clk);
#1;data_in = testData6[8340];
@(posedge clk);
#1;data_in = testData6[8341];
@(posedge clk);
#1;data_in = testData6[8342];
@(posedge clk);
#1;data_in = testData6[8343];
@(posedge clk);
#1;data_in = testData6[8344];
@(posedge clk);
#1;data_in = testData6[8345];
@(posedge clk);
#1;data_in = testData6[8346];
@(posedge clk);
#1;data_in = testData6[8347];
@(posedge clk);
#1;data_in = testData6[8348];
@(posedge clk);
#1;data_in = testData6[8349];
@(posedge clk);
#1;data_in = testData6[8350];
@(posedge clk);
#1;data_in = testData6[8351];
@(posedge clk);
#1;data_in = testData6[8352];
@(posedge clk);
#1;data_in = testData6[8353];
@(posedge clk);
#1;data_in = testData6[8354];
@(posedge clk);
#1;data_in = testData6[8355];
@(posedge clk);
#1;data_in = testData6[8356];
@(posedge clk);
#1;data_in = testData6[8357];
@(posedge clk);
#1;data_in = testData6[8358];
@(posedge clk);
#1;data_in = testData6[8359];
@(posedge clk);
#1;data_in = testData6[8360];
@(posedge clk);
#1;data_in = testData6[8361];
@(posedge clk);
#1;data_in = testData6[8362];
@(posedge clk);
#1;data_in = testData6[8363];
@(posedge clk);
#1;data_in = testData6[8364];
@(posedge clk);
#1;data_in = testData6[8365];
@(posedge clk);
#1;data_in = testData6[8366];
@(posedge clk);
#1;data_in = testData6[8367];
@(posedge clk);
#1;data_in = testData6[8368];
@(posedge clk);
#1;data_in = testData6[8369];
@(posedge clk);
#1;data_in = testData6[8370];
@(posedge clk);
#1;data_in = testData6[8371];
@(posedge clk);
#1;data_in = testData6[8372];
@(posedge clk);
#1;data_in = testData6[8373];
@(posedge clk);
#1;data_in = testData6[8374];
@(posedge clk);
#1;data_in = testData6[8375];
@(posedge clk);
#1;data_in = testData6[8376];
@(posedge clk);
#1;data_in = testData6[8377];
@(posedge clk);
#1;data_in = testData6[8378];
@(posedge clk);
#1;data_in = testData6[8379];
@(posedge clk);
#1;data_in = testData6[8380];
@(posedge clk);
#1;data_in = testData6[8381];
@(posedge clk);
#1;data_in = testData6[8382];
@(posedge clk);
#1;data_in = testData6[8383];
@(posedge clk);
#1;data_in = testData6[8384];
@(posedge clk);
#1;data_in = testData6[8385];
@(posedge clk);
#1;data_in = testData6[8386];
@(posedge clk);
#1;data_in = testData6[8387];
@(posedge clk);
#1;data_in = testData6[8388];
@(posedge clk);
#1;data_in = testData6[8389];
@(posedge clk);
#1;data_in = testData6[8390];
@(posedge clk);
#1;data_in = testData6[8391];
@(posedge clk);
#1;data_in = testData6[8392];
@(posedge clk);
#1;data_in = testData6[8393];
@(posedge clk);
#1;data_in = testData6[8394];
@(posedge clk);
#1;data_in = testData6[8395];
@(posedge clk);
#1;data_in = testData6[8396];
@(posedge clk);
#1;data_in = testData6[8397];
@(posedge clk);
#1;data_in = testData6[8398];
@(posedge clk);
#1;data_in = testData6[8399];
@(posedge clk);
#1;data_in = testData6[8400];
@(posedge clk);
#1;data_in = testData6[8401];
@(posedge clk);
#1;data_in = testData6[8402];
@(posedge clk);
#1;data_in = testData6[8403];
@(posedge clk);
#1;data_in = testData6[8404];
@(posedge clk);
#1;data_in = testData6[8405];
@(posedge clk);
#1;data_in = testData6[8406];
@(posedge clk);
#1;data_in = testData6[8407];
@(posedge clk);
#1;data_in = testData6[8408];
@(posedge clk);
#1;data_in = testData6[8409];
@(posedge clk);
#1;data_in = testData6[8410];
@(posedge clk);
#1;data_in = testData6[8411];
@(posedge clk);
#1;data_in = testData6[8412];
@(posedge clk);
#1;data_in = testData6[8413];
@(posedge clk);
#1;data_in = testData6[8414];
@(posedge clk);
#1;data_in = testData6[8415];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[8416]; 
@(posedge clk);
#1;data_in = testData6[8417];
@(posedge clk);
#1;data_in = testData6[8418];
@(posedge clk);
#1;data_in = testData6[8419];
@(posedge clk);
#1;data_in = testData6[8420];
@(posedge clk);
#1;data_in = testData6[8421];
@(posedge clk);
#1;data_in = testData6[8422];
@(posedge clk);
#1;data_in = testData6[8423];
@(posedge clk);
#1;data_in = testData6[8424];
@(posedge clk);
#1;data_in = testData6[8425];
@(posedge clk);
#1;data_in = testData6[8426];
@(posedge clk);
#1;data_in = testData6[8427];
@(posedge clk);
#1;data_in = testData6[8428];
@(posedge clk);
#1;data_in = testData6[8429];
@(posedge clk);
#1;data_in = testData6[8430];
@(posedge clk);
#1;data_in = testData6[8431];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[8432];
@(posedge clk);
#1;data_in = testData6[8433];
@(posedge clk);
#1;data_in = testData6[8434];
@(posedge clk);
#1;data_in = testData6[8435];
@(posedge clk);
#1;data_in = testData6[8436];
@(posedge clk);
#1;data_in = testData6[8437];
@(posedge clk);
#1;data_in = testData6[8438];
@(posedge clk);
#1;data_in = testData6[8439];
@(posedge clk);
#1;data_in = testData6[8440];
@(posedge clk);
#1;data_in = testData6[8441];
@(posedge clk);
#1;data_in = testData6[8442];
@(posedge clk);
#1;data_in = testData6[8443];
@(posedge clk);
#1;data_in = testData6[8444];
@(posedge clk);
#1;data_in = testData6[8445];
@(posedge clk);
#1;data_in = testData6[8446];
@(posedge clk);
#1;data_in = testData6[8447];
@(posedge clk);
#1;data_in = testData6[8448];
@(posedge clk);
#1;data_in = testData6[8449];
@(posedge clk);
#1;data_in = testData6[8450];
@(posedge clk);
#1;data_in = testData6[8451];
@(posedge clk);
#1;data_in = testData6[8452];
@(posedge clk);
#1;data_in = testData6[8453];
@(posedge clk);
#1;data_in = testData6[8454];
@(posedge clk);
#1;data_in = testData6[8455];
@(posedge clk);
#1;data_in = testData6[8456];
@(posedge clk);
#1;data_in = testData6[8457];
@(posedge clk);
#1;data_in = testData6[8458];
@(posedge clk);
#1;data_in = testData6[8459];
@(posedge clk);
#1;data_in = testData6[8460];
@(posedge clk);
#1;data_in = testData6[8461];
@(posedge clk);
#1;data_in = testData6[8462];
@(posedge clk);
#1;data_in = testData6[8463];
@(posedge clk);
#1;data_in = testData6[8464];
@(posedge clk);
#1;data_in = testData6[8465];
@(posedge clk);
#1;data_in = testData6[8466];
@(posedge clk);
#1;data_in = testData6[8467];
@(posedge clk);
#1;data_in = testData6[8468];
@(posedge clk);
#1;data_in = testData6[8469];
@(posedge clk);
#1;data_in = testData6[8470];
@(posedge clk);
#1;data_in = testData6[8471];
@(posedge clk);
#1;data_in = testData6[8472];
@(posedge clk);
#1;data_in = testData6[8473];
@(posedge clk);
#1;data_in = testData6[8474];
@(posedge clk);
#1;data_in = testData6[8475];
@(posedge clk);
#1;data_in = testData6[8476];
@(posedge clk);
#1;data_in = testData6[8477];
@(posedge clk);
#1;data_in = testData6[8478];
@(posedge clk);
#1;data_in = testData6[8479];
@(posedge clk);
#1;data_in = testData6[8480];
@(posedge clk);
#1;data_in = testData6[8481];
@(posedge clk);
#1;data_in = testData6[8482];
@(posedge clk);
#1;data_in = testData6[8483];
@(posedge clk);
#1;data_in = testData6[8484];
@(posedge clk);
#1;data_in = testData6[8485];
@(posedge clk);
#1;data_in = testData6[8486];
@(posedge clk);
#1;data_in = testData6[8487];
@(posedge clk);
#1;data_in = testData6[8488];
@(posedge clk);
#1;data_in = testData6[8489];
@(posedge clk);
#1;data_in = testData6[8490];
@(posedge clk);
#1;data_in = testData6[8491];
@(posedge clk);
#1;data_in = testData6[8492];
@(posedge clk);
#1;data_in = testData6[8493];
@(posedge clk);
#1;data_in = testData6[8494];
@(posedge clk);
#1;data_in = testData6[8495];
@(posedge clk);
#1;data_in = testData6[8496];
@(posedge clk);
#1;data_in = testData6[8497];
@(posedge clk);
#1;data_in = testData6[8498];
@(posedge clk);
#1;data_in = testData6[8499];
@(posedge clk);
#1;data_in = testData6[8500];
@(posedge clk);
#1;data_in = testData6[8501];
@(posedge clk);
#1;data_in = testData6[8502];
@(posedge clk);
#1;data_in = testData6[8503];
@(posedge clk);
#1;data_in = testData6[8504];
@(posedge clk);
#1;data_in = testData6[8505];
@(posedge clk);
#1;data_in = testData6[8506];
@(posedge clk);
#1;data_in = testData6[8507];
@(posedge clk);
#1;data_in = testData6[8508];
@(posedge clk);
#1;data_in = testData6[8509];
@(posedge clk);
#1;data_in = testData6[8510];
@(posedge clk);
#1;data_in = testData6[8511];
@(posedge clk);
#1;data_in = testData6[8512];
@(posedge clk);
#1;data_in = testData6[8513];
@(posedge clk);
#1;data_in = testData6[8514];
@(posedge clk);
#1;data_in = testData6[8515];
@(posedge clk);
#1;data_in = testData6[8516];
@(posedge clk);
#1;data_in = testData6[8517];
@(posedge clk);
#1;data_in = testData6[8518];
@(posedge clk);
#1;data_in = testData6[8519];
@(posedge clk);
#1;data_in = testData6[8520];
@(posedge clk);
#1;data_in = testData6[8521];
@(posedge clk);
#1;data_in = testData6[8522];
@(posedge clk);
#1;data_in = testData6[8523];
@(posedge clk);
#1;data_in = testData6[8524];
@(posedge clk);
#1;data_in = testData6[8525];
@(posedge clk);
#1;data_in = testData6[8526];
@(posedge clk);
#1;data_in = testData6[8527];
@(posedge clk);
#1;data_in = testData6[8528];
@(posedge clk);
#1;data_in = testData6[8529];
@(posedge clk);
#1;data_in = testData6[8530];
@(posedge clk);
#1;data_in = testData6[8531];
@(posedge clk);
#1;data_in = testData6[8532];
@(posedge clk);
#1;data_in = testData6[8533];
@(posedge clk);
#1;data_in = testData6[8534];
@(posedge clk);
#1;data_in = testData6[8535];
@(posedge clk);
#1;data_in = testData6[8536];
@(posedge clk);
#1;data_in = testData6[8537];
@(posedge clk);
#1;data_in = testData6[8538];
@(posedge clk);
#1;data_in = testData6[8539];
@(posedge clk);
#1;data_in = testData6[8540];
@(posedge clk);
#1;data_in = testData6[8541];
@(posedge clk);
#1;data_in = testData6[8542];
@(posedge clk);
#1;data_in = testData6[8543];
@(posedge clk);
#1;data_in = testData6[8544];
@(posedge clk);
#1;data_in = testData6[8545];
@(posedge clk);
#1;data_in = testData6[8546];
@(posedge clk);
#1;data_in = testData6[8547];
@(posedge clk);
#1;data_in = testData6[8548];
@(posedge clk);
#1;data_in = testData6[8549];
@(posedge clk);
#1;data_in = testData6[8550];
@(posedge clk);
#1;data_in = testData6[8551];
@(posedge clk);
#1;data_in = testData6[8552];
@(posedge clk);
#1;data_in = testData6[8553];
@(posedge clk);
#1;data_in = testData6[8554];
@(posedge clk);
#1;data_in = testData6[8555];
@(posedge clk);
#1;data_in = testData6[8556];
@(posedge clk);
#1;data_in = testData6[8557];
@(posedge clk);
#1;data_in = testData6[8558];
@(posedge clk);
#1;data_in = testData6[8559];
@(posedge clk);
#1;data_in = testData6[8560];
@(posedge clk);
#1;data_in = testData6[8561];
@(posedge clk);
#1;data_in = testData6[8562];
@(posedge clk);
#1;data_in = testData6[8563];
@(posedge clk);
#1;data_in = testData6[8564];
@(posedge clk);
#1;data_in = testData6[8565];
@(posedge clk);
#1;data_in = testData6[8566];
@(posedge clk);
#1;data_in = testData6[8567];
@(posedge clk);
#1;data_in = testData6[8568];
@(posedge clk);
#1;data_in = testData6[8569];
@(posedge clk);
#1;data_in = testData6[8570];
@(posedge clk);
#1;data_in = testData6[8571];
@(posedge clk);
#1;data_in = testData6[8572];
@(posedge clk);
#1;data_in = testData6[8573];
@(posedge clk);
#1;data_in = testData6[8574];
@(posedge clk);
#1;data_in = testData6[8575];
@(posedge clk);
#1;data_in = testData6[8576];
@(posedge clk);
#1;data_in = testData6[8577];
@(posedge clk);
#1;data_in = testData6[8578];
@(posedge clk);
#1;data_in = testData6[8579];
@(posedge clk);
#1;data_in = testData6[8580];
@(posedge clk);
#1;data_in = testData6[8581];
@(posedge clk);
#1;data_in = testData6[8582];
@(posedge clk);
#1;data_in = testData6[8583];
@(posedge clk);
#1;data_in = testData6[8584];
@(posedge clk);
#1;data_in = testData6[8585];
@(posedge clk);
#1;data_in = testData6[8586];
@(posedge clk);
#1;data_in = testData6[8587];
@(posedge clk);
#1;data_in = testData6[8588];
@(posedge clk);
#1;data_in = testData6[8589];
@(posedge clk);
#1;data_in = testData6[8590];
@(posedge clk);
#1;data_in = testData6[8591];
@(posedge clk);
#1;data_in = testData6[8592];
@(posedge clk);
#1;data_in = testData6[8593];
@(posedge clk);
#1;data_in = testData6[8594];
@(posedge clk);
#1;data_in = testData6[8595];
@(posedge clk);
#1;data_in = testData6[8596];
@(posedge clk);
#1;data_in = testData6[8597];
@(posedge clk);
#1;data_in = testData6[8598];
@(posedge clk);
#1;data_in = testData6[8599];
@(posedge clk);
#1;data_in = testData6[8600];
@(posedge clk);
#1;data_in = testData6[8601];
@(posedge clk);
#1;data_in = testData6[8602];
@(posedge clk);
#1;data_in = testData6[8603];
@(posedge clk);
#1;data_in = testData6[8604];
@(posedge clk);
#1;data_in = testData6[8605];
@(posedge clk);
#1;data_in = testData6[8606];
@(posedge clk);
#1;data_in = testData6[8607];
@(posedge clk);
#1;data_in = testData6[8608];
@(posedge clk);
#1;data_in = testData6[8609];
@(posedge clk);
#1;data_in = testData6[8610];
@(posedge clk);
#1;data_in = testData6[8611];
@(posedge clk);
#1;data_in = testData6[8612];
@(posedge clk);
#1;data_in = testData6[8613];
@(posedge clk);
#1;data_in = testData6[8614];
@(posedge clk);
#1;data_in = testData6[8615];
@(posedge clk);
#1;data_in = testData6[8616];
@(posedge clk);
#1;data_in = testData6[8617];
@(posedge clk);
#1;data_in = testData6[8618];
@(posedge clk);
#1;data_in = testData6[8619];
@(posedge clk);
#1;data_in = testData6[8620];
@(posedge clk);
#1;data_in = testData6[8621];
@(posedge clk);
#1;data_in = testData6[8622];
@(posedge clk);
#1;data_in = testData6[8623];
@(posedge clk);
#1;data_in = testData6[8624];
@(posedge clk);
#1;data_in = testData6[8625];
@(posedge clk);
#1;data_in = testData6[8626];
@(posedge clk);
#1;data_in = testData6[8627];
@(posedge clk);
#1;data_in = testData6[8628];
@(posedge clk);
#1;data_in = testData6[8629];
@(posedge clk);
#1;data_in = testData6[8630];
@(posedge clk);
#1;data_in = testData6[8631];
@(posedge clk);
#1;data_in = testData6[8632];
@(posedge clk);
#1;data_in = testData6[8633];
@(posedge clk);
#1;data_in = testData6[8634];
@(posedge clk);
#1;data_in = testData6[8635];
@(posedge clk);
#1;data_in = testData6[8636];
@(posedge clk);
#1;data_in = testData6[8637];
@(posedge clk);
#1;data_in = testData6[8638];
@(posedge clk);
#1;data_in = testData6[8639];
@(posedge clk);
#1;data_in = testData6[8640];
@(posedge clk);
#1;data_in = testData6[8641];
@(posedge clk);
#1;data_in = testData6[8642];
@(posedge clk);
#1;data_in = testData6[8643];
@(posedge clk);
#1;data_in = testData6[8644];
@(posedge clk);
#1;data_in = testData6[8645];
@(posedge clk);
#1;data_in = testData6[8646];
@(posedge clk);
#1;data_in = testData6[8647];
@(posedge clk);
#1;data_in = testData6[8648];
@(posedge clk);
#1;data_in = testData6[8649];
@(posedge clk);
#1;data_in = testData6[8650];
@(posedge clk);
#1;data_in = testData6[8651];
@(posedge clk);
#1;data_in = testData6[8652];
@(posedge clk);
#1;data_in = testData6[8653];
@(posedge clk);
#1;data_in = testData6[8654];
@(posedge clk);
#1;data_in = testData6[8655];
@(posedge clk);
#1;data_in = testData6[8656];
@(posedge clk);
#1;data_in = testData6[8657];
@(posedge clk);
#1;data_in = testData6[8658];
@(posedge clk);
#1;data_in = testData6[8659];
@(posedge clk);
#1;data_in = testData6[8660];
@(posedge clk);
#1;data_in = testData6[8661];
@(posedge clk);
#1;data_in = testData6[8662];
@(posedge clk);
#1;data_in = testData6[8663];
@(posedge clk);
#1;data_in = testData6[8664];
@(posedge clk);
#1;data_in = testData6[8665];
@(posedge clk);
#1;data_in = testData6[8666];
@(posedge clk);
#1;data_in = testData6[8667];
@(posedge clk);
#1;data_in = testData6[8668];
@(posedge clk);
#1;data_in = testData6[8669];
@(posedge clk);
#1;data_in = testData6[8670];
@(posedge clk);
#1;data_in = testData6[8671];
@(posedge clk);
#1;data_in = testData6[8672];
@(posedge clk);
#1;data_in = testData6[8673];
@(posedge clk);
#1;data_in = testData6[8674];
@(posedge clk);
#1;data_in = testData6[8675];
@(posedge clk);
#1;data_in = testData6[8676];
@(posedge clk);
#1;data_in = testData6[8677];
@(posedge clk);
#1;data_in = testData6[8678];
@(posedge clk);
#1;data_in = testData6[8679];
@(posedge clk);
#1;data_in = testData6[8680];
@(posedge clk);
#1;data_in = testData6[8681];
@(posedge clk);
#1;data_in = testData6[8682];
@(posedge clk);
#1;data_in = testData6[8683];
@(posedge clk);
#1;data_in = testData6[8684];
@(posedge clk);
#1;data_in = testData6[8685];
@(posedge clk);
#1;data_in = testData6[8686];
@(posedge clk);
#1;data_in = testData6[8687];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[8688]; 
@(posedge clk);
#1;data_in = testData6[8689];
@(posedge clk);
#1;data_in = testData6[8690];
@(posedge clk);
#1;data_in = testData6[8691];
@(posedge clk);
#1;data_in = testData6[8692];
@(posedge clk);
#1;data_in = testData6[8693];
@(posedge clk);
#1;data_in = testData6[8694];
@(posedge clk);
#1;data_in = testData6[8695];
@(posedge clk);
#1;data_in = testData6[8696];
@(posedge clk);
#1;data_in = testData6[8697];
@(posedge clk);
#1;data_in = testData6[8698];
@(posedge clk);
#1;data_in = testData6[8699];
@(posedge clk);
#1;data_in = testData6[8700];
@(posedge clk);
#1;data_in = testData6[8701];
@(posedge clk);
#1;data_in = testData6[8702];
@(posedge clk);
#1;data_in = testData6[8703];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[8704];
@(posedge clk);
#1;data_in = testData6[8705];
@(posedge clk);
#1;data_in = testData6[8706];
@(posedge clk);
#1;data_in = testData6[8707];
@(posedge clk);
#1;data_in = testData6[8708];
@(posedge clk);
#1;data_in = testData6[8709];
@(posedge clk);
#1;data_in = testData6[8710];
@(posedge clk);
#1;data_in = testData6[8711];
@(posedge clk);
#1;data_in = testData6[8712];
@(posedge clk);
#1;data_in = testData6[8713];
@(posedge clk);
#1;data_in = testData6[8714];
@(posedge clk);
#1;data_in = testData6[8715];
@(posedge clk);
#1;data_in = testData6[8716];
@(posedge clk);
#1;data_in = testData6[8717];
@(posedge clk);
#1;data_in = testData6[8718];
@(posedge clk);
#1;data_in = testData6[8719];
@(posedge clk);
#1;data_in = testData6[8720];
@(posedge clk);
#1;data_in = testData6[8721];
@(posedge clk);
#1;data_in = testData6[8722];
@(posedge clk);
#1;data_in = testData6[8723];
@(posedge clk);
#1;data_in = testData6[8724];
@(posedge clk);
#1;data_in = testData6[8725];
@(posedge clk);
#1;data_in = testData6[8726];
@(posedge clk);
#1;data_in = testData6[8727];
@(posedge clk);
#1;data_in = testData6[8728];
@(posedge clk);
#1;data_in = testData6[8729];
@(posedge clk);
#1;data_in = testData6[8730];
@(posedge clk);
#1;data_in = testData6[8731];
@(posedge clk);
#1;data_in = testData6[8732];
@(posedge clk);
#1;data_in = testData6[8733];
@(posedge clk);
#1;data_in = testData6[8734];
@(posedge clk);
#1;data_in = testData6[8735];
@(posedge clk);
#1;data_in = testData6[8736];
@(posedge clk);
#1;data_in = testData6[8737];
@(posedge clk);
#1;data_in = testData6[8738];
@(posedge clk);
#1;data_in = testData6[8739];
@(posedge clk);
#1;data_in = testData6[8740];
@(posedge clk);
#1;data_in = testData6[8741];
@(posedge clk);
#1;data_in = testData6[8742];
@(posedge clk);
#1;data_in = testData6[8743];
@(posedge clk);
#1;data_in = testData6[8744];
@(posedge clk);
#1;data_in = testData6[8745];
@(posedge clk);
#1;data_in = testData6[8746];
@(posedge clk);
#1;data_in = testData6[8747];
@(posedge clk);
#1;data_in = testData6[8748];
@(posedge clk);
#1;data_in = testData6[8749];
@(posedge clk);
#1;data_in = testData6[8750];
@(posedge clk);
#1;data_in = testData6[8751];
@(posedge clk);
#1;data_in = testData6[8752];
@(posedge clk);
#1;data_in = testData6[8753];
@(posedge clk);
#1;data_in = testData6[8754];
@(posedge clk);
#1;data_in = testData6[8755];
@(posedge clk);
#1;data_in = testData6[8756];
@(posedge clk);
#1;data_in = testData6[8757];
@(posedge clk);
#1;data_in = testData6[8758];
@(posedge clk);
#1;data_in = testData6[8759];
@(posedge clk);
#1;data_in = testData6[8760];
@(posedge clk);
#1;data_in = testData6[8761];
@(posedge clk);
#1;data_in = testData6[8762];
@(posedge clk);
#1;data_in = testData6[8763];
@(posedge clk);
#1;data_in = testData6[8764];
@(posedge clk);
#1;data_in = testData6[8765];
@(posedge clk);
#1;data_in = testData6[8766];
@(posedge clk);
#1;data_in = testData6[8767];
@(posedge clk);
#1;data_in = testData6[8768];
@(posedge clk);
#1;data_in = testData6[8769];
@(posedge clk);
#1;data_in = testData6[8770];
@(posedge clk);
#1;data_in = testData6[8771];
@(posedge clk);
#1;data_in = testData6[8772];
@(posedge clk);
#1;data_in = testData6[8773];
@(posedge clk);
#1;data_in = testData6[8774];
@(posedge clk);
#1;data_in = testData6[8775];
@(posedge clk);
#1;data_in = testData6[8776];
@(posedge clk);
#1;data_in = testData6[8777];
@(posedge clk);
#1;data_in = testData6[8778];
@(posedge clk);
#1;data_in = testData6[8779];
@(posedge clk);
#1;data_in = testData6[8780];
@(posedge clk);
#1;data_in = testData6[8781];
@(posedge clk);
#1;data_in = testData6[8782];
@(posedge clk);
#1;data_in = testData6[8783];
@(posedge clk);
#1;data_in = testData6[8784];
@(posedge clk);
#1;data_in = testData6[8785];
@(posedge clk);
#1;data_in = testData6[8786];
@(posedge clk);
#1;data_in = testData6[8787];
@(posedge clk);
#1;data_in = testData6[8788];
@(posedge clk);
#1;data_in = testData6[8789];
@(posedge clk);
#1;data_in = testData6[8790];
@(posedge clk);
#1;data_in = testData6[8791];
@(posedge clk);
#1;data_in = testData6[8792];
@(posedge clk);
#1;data_in = testData6[8793];
@(posedge clk);
#1;data_in = testData6[8794];
@(posedge clk);
#1;data_in = testData6[8795];
@(posedge clk);
#1;data_in = testData6[8796];
@(posedge clk);
#1;data_in = testData6[8797];
@(posedge clk);
#1;data_in = testData6[8798];
@(posedge clk);
#1;data_in = testData6[8799];
@(posedge clk);
#1;data_in = testData6[8800];
@(posedge clk);
#1;data_in = testData6[8801];
@(posedge clk);
#1;data_in = testData6[8802];
@(posedge clk);
#1;data_in = testData6[8803];
@(posedge clk);
#1;data_in = testData6[8804];
@(posedge clk);
#1;data_in = testData6[8805];
@(posedge clk);
#1;data_in = testData6[8806];
@(posedge clk);
#1;data_in = testData6[8807];
@(posedge clk);
#1;data_in = testData6[8808];
@(posedge clk);
#1;data_in = testData6[8809];
@(posedge clk);
#1;data_in = testData6[8810];
@(posedge clk);
#1;data_in = testData6[8811];
@(posedge clk);
#1;data_in = testData6[8812];
@(posedge clk);
#1;data_in = testData6[8813];
@(posedge clk);
#1;data_in = testData6[8814];
@(posedge clk);
#1;data_in = testData6[8815];
@(posedge clk);
#1;data_in = testData6[8816];
@(posedge clk);
#1;data_in = testData6[8817];
@(posedge clk);
#1;data_in = testData6[8818];
@(posedge clk);
#1;data_in = testData6[8819];
@(posedge clk);
#1;data_in = testData6[8820];
@(posedge clk);
#1;data_in = testData6[8821];
@(posedge clk);
#1;data_in = testData6[8822];
@(posedge clk);
#1;data_in = testData6[8823];
@(posedge clk);
#1;data_in = testData6[8824];
@(posedge clk);
#1;data_in = testData6[8825];
@(posedge clk);
#1;data_in = testData6[8826];
@(posedge clk);
#1;data_in = testData6[8827];
@(posedge clk);
#1;data_in = testData6[8828];
@(posedge clk);
#1;data_in = testData6[8829];
@(posedge clk);
#1;data_in = testData6[8830];
@(posedge clk);
#1;data_in = testData6[8831];
@(posedge clk);
#1;data_in = testData6[8832];
@(posedge clk);
#1;data_in = testData6[8833];
@(posedge clk);
#1;data_in = testData6[8834];
@(posedge clk);
#1;data_in = testData6[8835];
@(posedge clk);
#1;data_in = testData6[8836];
@(posedge clk);
#1;data_in = testData6[8837];
@(posedge clk);
#1;data_in = testData6[8838];
@(posedge clk);
#1;data_in = testData6[8839];
@(posedge clk);
#1;data_in = testData6[8840];
@(posedge clk);
#1;data_in = testData6[8841];
@(posedge clk);
#1;data_in = testData6[8842];
@(posedge clk);
#1;data_in = testData6[8843];
@(posedge clk);
#1;data_in = testData6[8844];
@(posedge clk);
#1;data_in = testData6[8845];
@(posedge clk);
#1;data_in = testData6[8846];
@(posedge clk);
#1;data_in = testData6[8847];
@(posedge clk);
#1;data_in = testData6[8848];
@(posedge clk);
#1;data_in = testData6[8849];
@(posedge clk);
#1;data_in = testData6[8850];
@(posedge clk);
#1;data_in = testData6[8851];
@(posedge clk);
#1;data_in = testData6[8852];
@(posedge clk);
#1;data_in = testData6[8853];
@(posedge clk);
#1;data_in = testData6[8854];
@(posedge clk);
#1;data_in = testData6[8855];
@(posedge clk);
#1;data_in = testData6[8856];
@(posedge clk);
#1;data_in = testData6[8857];
@(posedge clk);
#1;data_in = testData6[8858];
@(posedge clk);
#1;data_in = testData6[8859];
@(posedge clk);
#1;data_in = testData6[8860];
@(posedge clk);
#1;data_in = testData6[8861];
@(posedge clk);
#1;data_in = testData6[8862];
@(posedge clk);
#1;data_in = testData6[8863];
@(posedge clk);
#1;data_in = testData6[8864];
@(posedge clk);
#1;data_in = testData6[8865];
@(posedge clk);
#1;data_in = testData6[8866];
@(posedge clk);
#1;data_in = testData6[8867];
@(posedge clk);
#1;data_in = testData6[8868];
@(posedge clk);
#1;data_in = testData6[8869];
@(posedge clk);
#1;data_in = testData6[8870];
@(posedge clk);
#1;data_in = testData6[8871];
@(posedge clk);
#1;data_in = testData6[8872];
@(posedge clk);
#1;data_in = testData6[8873];
@(posedge clk);
#1;data_in = testData6[8874];
@(posedge clk);
#1;data_in = testData6[8875];
@(posedge clk);
#1;data_in = testData6[8876];
@(posedge clk);
#1;data_in = testData6[8877];
@(posedge clk);
#1;data_in = testData6[8878];
@(posedge clk);
#1;data_in = testData6[8879];
@(posedge clk);
#1;data_in = testData6[8880];
@(posedge clk);
#1;data_in = testData6[8881];
@(posedge clk);
#1;data_in = testData6[8882];
@(posedge clk);
#1;data_in = testData6[8883];
@(posedge clk);
#1;data_in = testData6[8884];
@(posedge clk);
#1;data_in = testData6[8885];
@(posedge clk);
#1;data_in = testData6[8886];
@(posedge clk);
#1;data_in = testData6[8887];
@(posedge clk);
#1;data_in = testData6[8888];
@(posedge clk);
#1;data_in = testData6[8889];
@(posedge clk);
#1;data_in = testData6[8890];
@(posedge clk);
#1;data_in = testData6[8891];
@(posedge clk);
#1;data_in = testData6[8892];
@(posedge clk);
#1;data_in = testData6[8893];
@(posedge clk);
#1;data_in = testData6[8894];
@(posedge clk);
#1;data_in = testData6[8895];
@(posedge clk);
#1;data_in = testData6[8896];
@(posedge clk);
#1;data_in = testData6[8897];
@(posedge clk);
#1;data_in = testData6[8898];
@(posedge clk);
#1;data_in = testData6[8899];
@(posedge clk);
#1;data_in = testData6[8900];
@(posedge clk);
#1;data_in = testData6[8901];
@(posedge clk);
#1;data_in = testData6[8902];
@(posedge clk);
#1;data_in = testData6[8903];
@(posedge clk);
#1;data_in = testData6[8904];
@(posedge clk);
#1;data_in = testData6[8905];
@(posedge clk);
#1;data_in = testData6[8906];
@(posedge clk);
#1;data_in = testData6[8907];
@(posedge clk);
#1;data_in = testData6[8908];
@(posedge clk);
#1;data_in = testData6[8909];
@(posedge clk);
#1;data_in = testData6[8910];
@(posedge clk);
#1;data_in = testData6[8911];
@(posedge clk);
#1;data_in = testData6[8912];
@(posedge clk);
#1;data_in = testData6[8913];
@(posedge clk);
#1;data_in = testData6[8914];
@(posedge clk);
#1;data_in = testData6[8915];
@(posedge clk);
#1;data_in = testData6[8916];
@(posedge clk);
#1;data_in = testData6[8917];
@(posedge clk);
#1;data_in = testData6[8918];
@(posedge clk);
#1;data_in = testData6[8919];
@(posedge clk);
#1;data_in = testData6[8920];
@(posedge clk);
#1;data_in = testData6[8921];
@(posedge clk);
#1;data_in = testData6[8922];
@(posedge clk);
#1;data_in = testData6[8923];
@(posedge clk);
#1;data_in = testData6[8924];
@(posedge clk);
#1;data_in = testData6[8925];
@(posedge clk);
#1;data_in = testData6[8926];
@(posedge clk);
#1;data_in = testData6[8927];
@(posedge clk);
#1;data_in = testData6[8928];
@(posedge clk);
#1;data_in = testData6[8929];
@(posedge clk);
#1;data_in = testData6[8930];
@(posedge clk);
#1;data_in = testData6[8931];
@(posedge clk);
#1;data_in = testData6[8932];
@(posedge clk);
#1;data_in = testData6[8933];
@(posedge clk);
#1;data_in = testData6[8934];
@(posedge clk);
#1;data_in = testData6[8935];
@(posedge clk);
#1;data_in = testData6[8936];
@(posedge clk);
#1;data_in = testData6[8937];
@(posedge clk);
#1;data_in = testData6[8938];
@(posedge clk);
#1;data_in = testData6[8939];
@(posedge clk);
#1;data_in = testData6[8940];
@(posedge clk);
#1;data_in = testData6[8941];
@(posedge clk);
#1;data_in = testData6[8942];
@(posedge clk);
#1;data_in = testData6[8943];
@(posedge clk);
#1;data_in = testData6[8944];
@(posedge clk);
#1;data_in = testData6[8945];
@(posedge clk);
#1;data_in = testData6[8946];
@(posedge clk);
#1;data_in = testData6[8947];
@(posedge clk);
#1;data_in = testData6[8948];
@(posedge clk);
#1;data_in = testData6[8949];
@(posedge clk);
#1;data_in = testData6[8950];
@(posedge clk);
#1;data_in = testData6[8951];
@(posedge clk);
#1;data_in = testData6[8952];
@(posedge clk);
#1;data_in = testData6[8953];
@(posedge clk);
#1;data_in = testData6[8954];
@(posedge clk);
#1;data_in = testData6[8955];
@(posedge clk);
#1;data_in = testData6[8956];
@(posedge clk);
#1;data_in = testData6[8957];
@(posedge clk);
#1;data_in = testData6[8958];
@(posedge clk);
#1;data_in = testData6[8959];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[8960]; 
@(posedge clk);
#1;data_in = testData6[8961];
@(posedge clk);
#1;data_in = testData6[8962];
@(posedge clk);
#1;data_in = testData6[8963];
@(posedge clk);
#1;data_in = testData6[8964];
@(posedge clk);
#1;data_in = testData6[8965];
@(posedge clk);
#1;data_in = testData6[8966];
@(posedge clk);
#1;data_in = testData6[8967];
@(posedge clk);
#1;data_in = testData6[8968];
@(posedge clk);
#1;data_in = testData6[8969];
@(posedge clk);
#1;data_in = testData6[8970];
@(posedge clk);
#1;data_in = testData6[8971];
@(posedge clk);
#1;data_in = testData6[8972];
@(posedge clk);
#1;data_in = testData6[8973];
@(posedge clk);
#1;data_in = testData6[8974];
@(posedge clk);
#1;data_in = testData6[8975];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[8976];
@(posedge clk);
#1;data_in = testData6[8977];
@(posedge clk);
#1;data_in = testData6[8978];
@(posedge clk);
#1;data_in = testData6[8979];
@(posedge clk);
#1;data_in = testData6[8980];
@(posedge clk);
#1;data_in = testData6[8981];
@(posedge clk);
#1;data_in = testData6[8982];
@(posedge clk);
#1;data_in = testData6[8983];
@(posedge clk);
#1;data_in = testData6[8984];
@(posedge clk);
#1;data_in = testData6[8985];
@(posedge clk);
#1;data_in = testData6[8986];
@(posedge clk);
#1;data_in = testData6[8987];
@(posedge clk);
#1;data_in = testData6[8988];
@(posedge clk);
#1;data_in = testData6[8989];
@(posedge clk);
#1;data_in = testData6[8990];
@(posedge clk);
#1;data_in = testData6[8991];
@(posedge clk);
#1;data_in = testData6[8992];
@(posedge clk);
#1;data_in = testData6[8993];
@(posedge clk);
#1;data_in = testData6[8994];
@(posedge clk);
#1;data_in = testData6[8995];
@(posedge clk);
#1;data_in = testData6[8996];
@(posedge clk);
#1;data_in = testData6[8997];
@(posedge clk);
#1;data_in = testData6[8998];
@(posedge clk);
#1;data_in = testData6[8999];
@(posedge clk);
#1;data_in = testData6[9000];
@(posedge clk);
#1;data_in = testData6[9001];
@(posedge clk);
#1;data_in = testData6[9002];
@(posedge clk);
#1;data_in = testData6[9003];
@(posedge clk);
#1;data_in = testData6[9004];
@(posedge clk);
#1;data_in = testData6[9005];
@(posedge clk);
#1;data_in = testData6[9006];
@(posedge clk);
#1;data_in = testData6[9007];
@(posedge clk);
#1;data_in = testData6[9008];
@(posedge clk);
#1;data_in = testData6[9009];
@(posedge clk);
#1;data_in = testData6[9010];
@(posedge clk);
#1;data_in = testData6[9011];
@(posedge clk);
#1;data_in = testData6[9012];
@(posedge clk);
#1;data_in = testData6[9013];
@(posedge clk);
#1;data_in = testData6[9014];
@(posedge clk);
#1;data_in = testData6[9015];
@(posedge clk);
#1;data_in = testData6[9016];
@(posedge clk);
#1;data_in = testData6[9017];
@(posedge clk);
#1;data_in = testData6[9018];
@(posedge clk);
#1;data_in = testData6[9019];
@(posedge clk);
#1;data_in = testData6[9020];
@(posedge clk);
#1;data_in = testData6[9021];
@(posedge clk);
#1;data_in = testData6[9022];
@(posedge clk);
#1;data_in = testData6[9023];
@(posedge clk);
#1;data_in = testData6[9024];
@(posedge clk);
#1;data_in = testData6[9025];
@(posedge clk);
#1;data_in = testData6[9026];
@(posedge clk);
#1;data_in = testData6[9027];
@(posedge clk);
#1;data_in = testData6[9028];
@(posedge clk);
#1;data_in = testData6[9029];
@(posedge clk);
#1;data_in = testData6[9030];
@(posedge clk);
#1;data_in = testData6[9031];
@(posedge clk);
#1;data_in = testData6[9032];
@(posedge clk);
#1;data_in = testData6[9033];
@(posedge clk);
#1;data_in = testData6[9034];
@(posedge clk);
#1;data_in = testData6[9035];
@(posedge clk);
#1;data_in = testData6[9036];
@(posedge clk);
#1;data_in = testData6[9037];
@(posedge clk);
#1;data_in = testData6[9038];
@(posedge clk);
#1;data_in = testData6[9039];
@(posedge clk);
#1;data_in = testData6[9040];
@(posedge clk);
#1;data_in = testData6[9041];
@(posedge clk);
#1;data_in = testData6[9042];
@(posedge clk);
#1;data_in = testData6[9043];
@(posedge clk);
#1;data_in = testData6[9044];
@(posedge clk);
#1;data_in = testData6[9045];
@(posedge clk);
#1;data_in = testData6[9046];
@(posedge clk);
#1;data_in = testData6[9047];
@(posedge clk);
#1;data_in = testData6[9048];
@(posedge clk);
#1;data_in = testData6[9049];
@(posedge clk);
#1;data_in = testData6[9050];
@(posedge clk);
#1;data_in = testData6[9051];
@(posedge clk);
#1;data_in = testData6[9052];
@(posedge clk);
#1;data_in = testData6[9053];
@(posedge clk);
#1;data_in = testData6[9054];
@(posedge clk);
#1;data_in = testData6[9055];
@(posedge clk);
#1;data_in = testData6[9056];
@(posedge clk);
#1;data_in = testData6[9057];
@(posedge clk);
#1;data_in = testData6[9058];
@(posedge clk);
#1;data_in = testData6[9059];
@(posedge clk);
#1;data_in = testData6[9060];
@(posedge clk);
#1;data_in = testData6[9061];
@(posedge clk);
#1;data_in = testData6[9062];
@(posedge clk);
#1;data_in = testData6[9063];
@(posedge clk);
#1;data_in = testData6[9064];
@(posedge clk);
#1;data_in = testData6[9065];
@(posedge clk);
#1;data_in = testData6[9066];
@(posedge clk);
#1;data_in = testData6[9067];
@(posedge clk);
#1;data_in = testData6[9068];
@(posedge clk);
#1;data_in = testData6[9069];
@(posedge clk);
#1;data_in = testData6[9070];
@(posedge clk);
#1;data_in = testData6[9071];
@(posedge clk);
#1;data_in = testData6[9072];
@(posedge clk);
#1;data_in = testData6[9073];
@(posedge clk);
#1;data_in = testData6[9074];
@(posedge clk);
#1;data_in = testData6[9075];
@(posedge clk);
#1;data_in = testData6[9076];
@(posedge clk);
#1;data_in = testData6[9077];
@(posedge clk);
#1;data_in = testData6[9078];
@(posedge clk);
#1;data_in = testData6[9079];
@(posedge clk);
#1;data_in = testData6[9080];
@(posedge clk);
#1;data_in = testData6[9081];
@(posedge clk);
#1;data_in = testData6[9082];
@(posedge clk);
#1;data_in = testData6[9083];
@(posedge clk);
#1;data_in = testData6[9084];
@(posedge clk);
#1;data_in = testData6[9085];
@(posedge clk);
#1;data_in = testData6[9086];
@(posedge clk);
#1;data_in = testData6[9087];
@(posedge clk);
#1;data_in = testData6[9088];
@(posedge clk);
#1;data_in = testData6[9089];
@(posedge clk);
#1;data_in = testData6[9090];
@(posedge clk);
#1;data_in = testData6[9091];
@(posedge clk);
#1;data_in = testData6[9092];
@(posedge clk);
#1;data_in = testData6[9093];
@(posedge clk);
#1;data_in = testData6[9094];
@(posedge clk);
#1;data_in = testData6[9095];
@(posedge clk);
#1;data_in = testData6[9096];
@(posedge clk);
#1;data_in = testData6[9097];
@(posedge clk);
#1;data_in = testData6[9098];
@(posedge clk);
#1;data_in = testData6[9099];
@(posedge clk);
#1;data_in = testData6[9100];
@(posedge clk);
#1;data_in = testData6[9101];
@(posedge clk);
#1;data_in = testData6[9102];
@(posedge clk);
#1;data_in = testData6[9103];
@(posedge clk);
#1;data_in = testData6[9104];
@(posedge clk);
#1;data_in = testData6[9105];
@(posedge clk);
#1;data_in = testData6[9106];
@(posedge clk);
#1;data_in = testData6[9107];
@(posedge clk);
#1;data_in = testData6[9108];
@(posedge clk);
#1;data_in = testData6[9109];
@(posedge clk);
#1;data_in = testData6[9110];
@(posedge clk);
#1;data_in = testData6[9111];
@(posedge clk);
#1;data_in = testData6[9112];
@(posedge clk);
#1;data_in = testData6[9113];
@(posedge clk);
#1;data_in = testData6[9114];
@(posedge clk);
#1;data_in = testData6[9115];
@(posedge clk);
#1;data_in = testData6[9116];
@(posedge clk);
#1;data_in = testData6[9117];
@(posedge clk);
#1;data_in = testData6[9118];
@(posedge clk);
#1;data_in = testData6[9119];
@(posedge clk);
#1;data_in = testData6[9120];
@(posedge clk);
#1;data_in = testData6[9121];
@(posedge clk);
#1;data_in = testData6[9122];
@(posedge clk);
#1;data_in = testData6[9123];
@(posedge clk);
#1;data_in = testData6[9124];
@(posedge clk);
#1;data_in = testData6[9125];
@(posedge clk);
#1;data_in = testData6[9126];
@(posedge clk);
#1;data_in = testData6[9127];
@(posedge clk);
#1;data_in = testData6[9128];
@(posedge clk);
#1;data_in = testData6[9129];
@(posedge clk);
#1;data_in = testData6[9130];
@(posedge clk);
#1;data_in = testData6[9131];
@(posedge clk);
#1;data_in = testData6[9132];
@(posedge clk);
#1;data_in = testData6[9133];
@(posedge clk);
#1;data_in = testData6[9134];
@(posedge clk);
#1;data_in = testData6[9135];
@(posedge clk);
#1;data_in = testData6[9136];
@(posedge clk);
#1;data_in = testData6[9137];
@(posedge clk);
#1;data_in = testData6[9138];
@(posedge clk);
#1;data_in = testData6[9139];
@(posedge clk);
#1;data_in = testData6[9140];
@(posedge clk);
#1;data_in = testData6[9141];
@(posedge clk);
#1;data_in = testData6[9142];
@(posedge clk);
#1;data_in = testData6[9143];
@(posedge clk);
#1;data_in = testData6[9144];
@(posedge clk);
#1;data_in = testData6[9145];
@(posedge clk);
#1;data_in = testData6[9146];
@(posedge clk);
#1;data_in = testData6[9147];
@(posedge clk);
#1;data_in = testData6[9148];
@(posedge clk);
#1;data_in = testData6[9149];
@(posedge clk);
#1;data_in = testData6[9150];
@(posedge clk);
#1;data_in = testData6[9151];
@(posedge clk);
#1;data_in = testData6[9152];
@(posedge clk);
#1;data_in = testData6[9153];
@(posedge clk);
#1;data_in = testData6[9154];
@(posedge clk);
#1;data_in = testData6[9155];
@(posedge clk);
#1;data_in = testData6[9156];
@(posedge clk);
#1;data_in = testData6[9157];
@(posedge clk);
#1;data_in = testData6[9158];
@(posedge clk);
#1;data_in = testData6[9159];
@(posedge clk);
#1;data_in = testData6[9160];
@(posedge clk);
#1;data_in = testData6[9161];
@(posedge clk);
#1;data_in = testData6[9162];
@(posedge clk);
#1;data_in = testData6[9163];
@(posedge clk);
#1;data_in = testData6[9164];
@(posedge clk);
#1;data_in = testData6[9165];
@(posedge clk);
#1;data_in = testData6[9166];
@(posedge clk);
#1;data_in = testData6[9167];
@(posedge clk);
#1;data_in = testData6[9168];
@(posedge clk);
#1;data_in = testData6[9169];
@(posedge clk);
#1;data_in = testData6[9170];
@(posedge clk);
#1;data_in = testData6[9171];
@(posedge clk);
#1;data_in = testData6[9172];
@(posedge clk);
#1;data_in = testData6[9173];
@(posedge clk);
#1;data_in = testData6[9174];
@(posedge clk);
#1;data_in = testData6[9175];
@(posedge clk);
#1;data_in = testData6[9176];
@(posedge clk);
#1;data_in = testData6[9177];
@(posedge clk);
#1;data_in = testData6[9178];
@(posedge clk);
#1;data_in = testData6[9179];
@(posedge clk);
#1;data_in = testData6[9180];
@(posedge clk);
#1;data_in = testData6[9181];
@(posedge clk);
#1;data_in = testData6[9182];
@(posedge clk);
#1;data_in = testData6[9183];
@(posedge clk);
#1;data_in = testData6[9184];
@(posedge clk);
#1;data_in = testData6[9185];
@(posedge clk);
#1;data_in = testData6[9186];
@(posedge clk);
#1;data_in = testData6[9187];
@(posedge clk);
#1;data_in = testData6[9188];
@(posedge clk);
#1;data_in = testData6[9189];
@(posedge clk);
#1;data_in = testData6[9190];
@(posedge clk);
#1;data_in = testData6[9191];
@(posedge clk);
#1;data_in = testData6[9192];
@(posedge clk);
#1;data_in = testData6[9193];
@(posedge clk);
#1;data_in = testData6[9194];
@(posedge clk);
#1;data_in = testData6[9195];
@(posedge clk);
#1;data_in = testData6[9196];
@(posedge clk);
#1;data_in = testData6[9197];
@(posedge clk);
#1;data_in = testData6[9198];
@(posedge clk);
#1;data_in = testData6[9199];
@(posedge clk);
#1;data_in = testData6[9200];
@(posedge clk);
#1;data_in = testData6[9201];
@(posedge clk);
#1;data_in = testData6[9202];
@(posedge clk);
#1;data_in = testData6[9203];
@(posedge clk);
#1;data_in = testData6[9204];
@(posedge clk);
#1;data_in = testData6[9205];
@(posedge clk);
#1;data_in = testData6[9206];
@(posedge clk);
#1;data_in = testData6[9207];
@(posedge clk);
#1;data_in = testData6[9208];
@(posedge clk);
#1;data_in = testData6[9209];
@(posedge clk);
#1;data_in = testData6[9210];
@(posedge clk);
#1;data_in = testData6[9211];
@(posedge clk);
#1;data_in = testData6[9212];
@(posedge clk);
#1;data_in = testData6[9213];
@(posedge clk);
#1;data_in = testData6[9214];
@(posedge clk);
#1;data_in = testData6[9215];
@(posedge clk);
#1;data_in = testData6[9216];
@(posedge clk);
#1;data_in = testData6[9217];
@(posedge clk);
#1;data_in = testData6[9218];
@(posedge clk);
#1;data_in = testData6[9219];
@(posedge clk);
#1;data_in = testData6[9220];
@(posedge clk);
#1;data_in = testData6[9221];
@(posedge clk);
#1;data_in = testData6[9222];
@(posedge clk);
#1;data_in = testData6[9223];
@(posedge clk);
#1;data_in = testData6[9224];
@(posedge clk);
#1;data_in = testData6[9225];
@(posedge clk);
#1;data_in = testData6[9226];
@(posedge clk);
#1;data_in = testData6[9227];
@(posedge clk);
#1;data_in = testData6[9228];
@(posedge clk);
#1;data_in = testData6[9229];
@(posedge clk);
#1;data_in = testData6[9230];
@(posedge clk);
#1;data_in = testData6[9231];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[9232]; 
@(posedge clk);
#1;data_in = testData6[9233];
@(posedge clk);
#1;data_in = testData6[9234];
@(posedge clk);
#1;data_in = testData6[9235];
@(posedge clk);
#1;data_in = testData6[9236];
@(posedge clk);
#1;data_in = testData6[9237];
@(posedge clk);
#1;data_in = testData6[9238];
@(posedge clk);
#1;data_in = testData6[9239];
@(posedge clk);
#1;data_in = testData6[9240];
@(posedge clk);
#1;data_in = testData6[9241];
@(posedge clk);
#1;data_in = testData6[9242];
@(posedge clk);
#1;data_in = testData6[9243];
@(posedge clk);
#1;data_in = testData6[9244];
@(posedge clk);
#1;data_in = testData6[9245];
@(posedge clk);
#1;data_in = testData6[9246];
@(posedge clk);
#1;data_in = testData6[9247];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[9248];
@(posedge clk);
#1;data_in = testData6[9249];
@(posedge clk);
#1;data_in = testData6[9250];
@(posedge clk);
#1;data_in = testData6[9251];
@(posedge clk);
#1;data_in = testData6[9252];
@(posedge clk);
#1;data_in = testData6[9253];
@(posedge clk);
#1;data_in = testData6[9254];
@(posedge clk);
#1;data_in = testData6[9255];
@(posedge clk);
#1;data_in = testData6[9256];
@(posedge clk);
#1;data_in = testData6[9257];
@(posedge clk);
#1;data_in = testData6[9258];
@(posedge clk);
#1;data_in = testData6[9259];
@(posedge clk);
#1;data_in = testData6[9260];
@(posedge clk);
#1;data_in = testData6[9261];
@(posedge clk);
#1;data_in = testData6[9262];
@(posedge clk);
#1;data_in = testData6[9263];
@(posedge clk);
#1;data_in = testData6[9264];
@(posedge clk);
#1;data_in = testData6[9265];
@(posedge clk);
#1;data_in = testData6[9266];
@(posedge clk);
#1;data_in = testData6[9267];
@(posedge clk);
#1;data_in = testData6[9268];
@(posedge clk);
#1;data_in = testData6[9269];
@(posedge clk);
#1;data_in = testData6[9270];
@(posedge clk);
#1;data_in = testData6[9271];
@(posedge clk);
#1;data_in = testData6[9272];
@(posedge clk);
#1;data_in = testData6[9273];
@(posedge clk);
#1;data_in = testData6[9274];
@(posedge clk);
#1;data_in = testData6[9275];
@(posedge clk);
#1;data_in = testData6[9276];
@(posedge clk);
#1;data_in = testData6[9277];
@(posedge clk);
#1;data_in = testData6[9278];
@(posedge clk);
#1;data_in = testData6[9279];
@(posedge clk);
#1;data_in = testData6[9280];
@(posedge clk);
#1;data_in = testData6[9281];
@(posedge clk);
#1;data_in = testData6[9282];
@(posedge clk);
#1;data_in = testData6[9283];
@(posedge clk);
#1;data_in = testData6[9284];
@(posedge clk);
#1;data_in = testData6[9285];
@(posedge clk);
#1;data_in = testData6[9286];
@(posedge clk);
#1;data_in = testData6[9287];
@(posedge clk);
#1;data_in = testData6[9288];
@(posedge clk);
#1;data_in = testData6[9289];
@(posedge clk);
#1;data_in = testData6[9290];
@(posedge clk);
#1;data_in = testData6[9291];
@(posedge clk);
#1;data_in = testData6[9292];
@(posedge clk);
#1;data_in = testData6[9293];
@(posedge clk);
#1;data_in = testData6[9294];
@(posedge clk);
#1;data_in = testData6[9295];
@(posedge clk);
#1;data_in = testData6[9296];
@(posedge clk);
#1;data_in = testData6[9297];
@(posedge clk);
#1;data_in = testData6[9298];
@(posedge clk);
#1;data_in = testData6[9299];
@(posedge clk);
#1;data_in = testData6[9300];
@(posedge clk);
#1;data_in = testData6[9301];
@(posedge clk);
#1;data_in = testData6[9302];
@(posedge clk);
#1;data_in = testData6[9303];
@(posedge clk);
#1;data_in = testData6[9304];
@(posedge clk);
#1;data_in = testData6[9305];
@(posedge clk);
#1;data_in = testData6[9306];
@(posedge clk);
#1;data_in = testData6[9307];
@(posedge clk);
#1;data_in = testData6[9308];
@(posedge clk);
#1;data_in = testData6[9309];
@(posedge clk);
#1;data_in = testData6[9310];
@(posedge clk);
#1;data_in = testData6[9311];
@(posedge clk);
#1;data_in = testData6[9312];
@(posedge clk);
#1;data_in = testData6[9313];
@(posedge clk);
#1;data_in = testData6[9314];
@(posedge clk);
#1;data_in = testData6[9315];
@(posedge clk);
#1;data_in = testData6[9316];
@(posedge clk);
#1;data_in = testData6[9317];
@(posedge clk);
#1;data_in = testData6[9318];
@(posedge clk);
#1;data_in = testData6[9319];
@(posedge clk);
#1;data_in = testData6[9320];
@(posedge clk);
#1;data_in = testData6[9321];
@(posedge clk);
#1;data_in = testData6[9322];
@(posedge clk);
#1;data_in = testData6[9323];
@(posedge clk);
#1;data_in = testData6[9324];
@(posedge clk);
#1;data_in = testData6[9325];
@(posedge clk);
#1;data_in = testData6[9326];
@(posedge clk);
#1;data_in = testData6[9327];
@(posedge clk);
#1;data_in = testData6[9328];
@(posedge clk);
#1;data_in = testData6[9329];
@(posedge clk);
#1;data_in = testData6[9330];
@(posedge clk);
#1;data_in = testData6[9331];
@(posedge clk);
#1;data_in = testData6[9332];
@(posedge clk);
#1;data_in = testData6[9333];
@(posedge clk);
#1;data_in = testData6[9334];
@(posedge clk);
#1;data_in = testData6[9335];
@(posedge clk);
#1;data_in = testData6[9336];
@(posedge clk);
#1;data_in = testData6[9337];
@(posedge clk);
#1;data_in = testData6[9338];
@(posedge clk);
#1;data_in = testData6[9339];
@(posedge clk);
#1;data_in = testData6[9340];
@(posedge clk);
#1;data_in = testData6[9341];
@(posedge clk);
#1;data_in = testData6[9342];
@(posedge clk);
#1;data_in = testData6[9343];
@(posedge clk);
#1;data_in = testData6[9344];
@(posedge clk);
#1;data_in = testData6[9345];
@(posedge clk);
#1;data_in = testData6[9346];
@(posedge clk);
#1;data_in = testData6[9347];
@(posedge clk);
#1;data_in = testData6[9348];
@(posedge clk);
#1;data_in = testData6[9349];
@(posedge clk);
#1;data_in = testData6[9350];
@(posedge clk);
#1;data_in = testData6[9351];
@(posedge clk);
#1;data_in = testData6[9352];
@(posedge clk);
#1;data_in = testData6[9353];
@(posedge clk);
#1;data_in = testData6[9354];
@(posedge clk);
#1;data_in = testData6[9355];
@(posedge clk);
#1;data_in = testData6[9356];
@(posedge clk);
#1;data_in = testData6[9357];
@(posedge clk);
#1;data_in = testData6[9358];
@(posedge clk);
#1;data_in = testData6[9359];
@(posedge clk);
#1;data_in = testData6[9360];
@(posedge clk);
#1;data_in = testData6[9361];
@(posedge clk);
#1;data_in = testData6[9362];
@(posedge clk);
#1;data_in = testData6[9363];
@(posedge clk);
#1;data_in = testData6[9364];
@(posedge clk);
#1;data_in = testData6[9365];
@(posedge clk);
#1;data_in = testData6[9366];
@(posedge clk);
#1;data_in = testData6[9367];
@(posedge clk);
#1;data_in = testData6[9368];
@(posedge clk);
#1;data_in = testData6[9369];
@(posedge clk);
#1;data_in = testData6[9370];
@(posedge clk);
#1;data_in = testData6[9371];
@(posedge clk);
#1;data_in = testData6[9372];
@(posedge clk);
#1;data_in = testData6[9373];
@(posedge clk);
#1;data_in = testData6[9374];
@(posedge clk);
#1;data_in = testData6[9375];
@(posedge clk);
#1;data_in = testData6[9376];
@(posedge clk);
#1;data_in = testData6[9377];
@(posedge clk);
#1;data_in = testData6[9378];
@(posedge clk);
#1;data_in = testData6[9379];
@(posedge clk);
#1;data_in = testData6[9380];
@(posedge clk);
#1;data_in = testData6[9381];
@(posedge clk);
#1;data_in = testData6[9382];
@(posedge clk);
#1;data_in = testData6[9383];
@(posedge clk);
#1;data_in = testData6[9384];
@(posedge clk);
#1;data_in = testData6[9385];
@(posedge clk);
#1;data_in = testData6[9386];
@(posedge clk);
#1;data_in = testData6[9387];
@(posedge clk);
#1;data_in = testData6[9388];
@(posedge clk);
#1;data_in = testData6[9389];
@(posedge clk);
#1;data_in = testData6[9390];
@(posedge clk);
#1;data_in = testData6[9391];
@(posedge clk);
#1;data_in = testData6[9392];
@(posedge clk);
#1;data_in = testData6[9393];
@(posedge clk);
#1;data_in = testData6[9394];
@(posedge clk);
#1;data_in = testData6[9395];
@(posedge clk);
#1;data_in = testData6[9396];
@(posedge clk);
#1;data_in = testData6[9397];
@(posedge clk);
#1;data_in = testData6[9398];
@(posedge clk);
#1;data_in = testData6[9399];
@(posedge clk);
#1;data_in = testData6[9400];
@(posedge clk);
#1;data_in = testData6[9401];
@(posedge clk);
#1;data_in = testData6[9402];
@(posedge clk);
#1;data_in = testData6[9403];
@(posedge clk);
#1;data_in = testData6[9404];
@(posedge clk);
#1;data_in = testData6[9405];
@(posedge clk);
#1;data_in = testData6[9406];
@(posedge clk);
#1;data_in = testData6[9407];
@(posedge clk);
#1;data_in = testData6[9408];
@(posedge clk);
#1;data_in = testData6[9409];
@(posedge clk);
#1;data_in = testData6[9410];
@(posedge clk);
#1;data_in = testData6[9411];
@(posedge clk);
#1;data_in = testData6[9412];
@(posedge clk);
#1;data_in = testData6[9413];
@(posedge clk);
#1;data_in = testData6[9414];
@(posedge clk);
#1;data_in = testData6[9415];
@(posedge clk);
#1;data_in = testData6[9416];
@(posedge clk);
#1;data_in = testData6[9417];
@(posedge clk);
#1;data_in = testData6[9418];
@(posedge clk);
#1;data_in = testData6[9419];
@(posedge clk);
#1;data_in = testData6[9420];
@(posedge clk);
#1;data_in = testData6[9421];
@(posedge clk);
#1;data_in = testData6[9422];
@(posedge clk);
#1;data_in = testData6[9423];
@(posedge clk);
#1;data_in = testData6[9424];
@(posedge clk);
#1;data_in = testData6[9425];
@(posedge clk);
#1;data_in = testData6[9426];
@(posedge clk);
#1;data_in = testData6[9427];
@(posedge clk);
#1;data_in = testData6[9428];
@(posedge clk);
#1;data_in = testData6[9429];
@(posedge clk);
#1;data_in = testData6[9430];
@(posedge clk);
#1;data_in = testData6[9431];
@(posedge clk);
#1;data_in = testData6[9432];
@(posedge clk);
#1;data_in = testData6[9433];
@(posedge clk);
#1;data_in = testData6[9434];
@(posedge clk);
#1;data_in = testData6[9435];
@(posedge clk);
#1;data_in = testData6[9436];
@(posedge clk);
#1;data_in = testData6[9437];
@(posedge clk);
#1;data_in = testData6[9438];
@(posedge clk);
#1;data_in = testData6[9439];
@(posedge clk);
#1;data_in = testData6[9440];
@(posedge clk);
#1;data_in = testData6[9441];
@(posedge clk);
#1;data_in = testData6[9442];
@(posedge clk);
#1;data_in = testData6[9443];
@(posedge clk);
#1;data_in = testData6[9444];
@(posedge clk);
#1;data_in = testData6[9445];
@(posedge clk);
#1;data_in = testData6[9446];
@(posedge clk);
#1;data_in = testData6[9447];
@(posedge clk);
#1;data_in = testData6[9448];
@(posedge clk);
#1;data_in = testData6[9449];
@(posedge clk);
#1;data_in = testData6[9450];
@(posedge clk);
#1;data_in = testData6[9451];
@(posedge clk);
#1;data_in = testData6[9452];
@(posedge clk);
#1;data_in = testData6[9453];
@(posedge clk);
#1;data_in = testData6[9454];
@(posedge clk);
#1;data_in = testData6[9455];
@(posedge clk);
#1;data_in = testData6[9456];
@(posedge clk);
#1;data_in = testData6[9457];
@(posedge clk);
#1;data_in = testData6[9458];
@(posedge clk);
#1;data_in = testData6[9459];
@(posedge clk);
#1;data_in = testData6[9460];
@(posedge clk);
#1;data_in = testData6[9461];
@(posedge clk);
#1;data_in = testData6[9462];
@(posedge clk);
#1;data_in = testData6[9463];
@(posedge clk);
#1;data_in = testData6[9464];
@(posedge clk);
#1;data_in = testData6[9465];
@(posedge clk);
#1;data_in = testData6[9466];
@(posedge clk);
#1;data_in = testData6[9467];
@(posedge clk);
#1;data_in = testData6[9468];
@(posedge clk);
#1;data_in = testData6[9469];
@(posedge clk);
#1;data_in = testData6[9470];
@(posedge clk);
#1;data_in = testData6[9471];
@(posedge clk);
#1;data_in = testData6[9472];
@(posedge clk);
#1;data_in = testData6[9473];
@(posedge clk);
#1;data_in = testData6[9474];
@(posedge clk);
#1;data_in = testData6[9475];
@(posedge clk);
#1;data_in = testData6[9476];
@(posedge clk);
#1;data_in = testData6[9477];
@(posedge clk);
#1;data_in = testData6[9478];
@(posedge clk);
#1;data_in = testData6[9479];
@(posedge clk);
#1;data_in = testData6[9480];
@(posedge clk);
#1;data_in = testData6[9481];
@(posedge clk);
#1;data_in = testData6[9482];
@(posedge clk);
#1;data_in = testData6[9483];
@(posedge clk);
#1;data_in = testData6[9484];
@(posedge clk);
#1;data_in = testData6[9485];
@(posedge clk);
#1;data_in = testData6[9486];
@(posedge clk);
#1;data_in = testData6[9487];
@(posedge clk);
#1;data_in = testData6[9488];
@(posedge clk);
#1;data_in = testData6[9489];
@(posedge clk);
#1;data_in = testData6[9490];
@(posedge clk);
#1;data_in = testData6[9491];
@(posedge clk);
#1;data_in = testData6[9492];
@(posedge clk);
#1;data_in = testData6[9493];
@(posedge clk);
#1;data_in = testData6[9494];
@(posedge clk);
#1;data_in = testData6[9495];
@(posedge clk);
#1;data_in = testData6[9496];
@(posedge clk);
#1;data_in = testData6[9497];
@(posedge clk);
#1;data_in = testData6[9498];
@(posedge clk);
#1;data_in = testData6[9499];
@(posedge clk);
#1;data_in = testData6[9500];
@(posedge clk);
#1;data_in = testData6[9501];
@(posedge clk);
#1;data_in = testData6[9502];
@(posedge clk);
#1;data_in = testData6[9503];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[9504]; 
@(posedge clk);
#1;data_in = testData6[9505];
@(posedge clk);
#1;data_in = testData6[9506];
@(posedge clk);
#1;data_in = testData6[9507];
@(posedge clk);
#1;data_in = testData6[9508];
@(posedge clk);
#1;data_in = testData6[9509];
@(posedge clk);
#1;data_in = testData6[9510];
@(posedge clk);
#1;data_in = testData6[9511];
@(posedge clk);
#1;data_in = testData6[9512];
@(posedge clk);
#1;data_in = testData6[9513];
@(posedge clk);
#1;data_in = testData6[9514];
@(posedge clk);
#1;data_in = testData6[9515];
@(posedge clk);
#1;data_in = testData6[9516];
@(posedge clk);
#1;data_in = testData6[9517];
@(posedge clk);
#1;data_in = testData6[9518];
@(posedge clk);
#1;data_in = testData6[9519];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[9520];
@(posedge clk);
#1;data_in = testData6[9521];
@(posedge clk);
#1;data_in = testData6[9522];
@(posedge clk);
#1;data_in = testData6[9523];
@(posedge clk);
#1;data_in = testData6[9524];
@(posedge clk);
#1;data_in = testData6[9525];
@(posedge clk);
#1;data_in = testData6[9526];
@(posedge clk);
#1;data_in = testData6[9527];
@(posedge clk);
#1;data_in = testData6[9528];
@(posedge clk);
#1;data_in = testData6[9529];
@(posedge clk);
#1;data_in = testData6[9530];
@(posedge clk);
#1;data_in = testData6[9531];
@(posedge clk);
#1;data_in = testData6[9532];
@(posedge clk);
#1;data_in = testData6[9533];
@(posedge clk);
#1;data_in = testData6[9534];
@(posedge clk);
#1;data_in = testData6[9535];
@(posedge clk);
#1;data_in = testData6[9536];
@(posedge clk);
#1;data_in = testData6[9537];
@(posedge clk);
#1;data_in = testData6[9538];
@(posedge clk);
#1;data_in = testData6[9539];
@(posedge clk);
#1;data_in = testData6[9540];
@(posedge clk);
#1;data_in = testData6[9541];
@(posedge clk);
#1;data_in = testData6[9542];
@(posedge clk);
#1;data_in = testData6[9543];
@(posedge clk);
#1;data_in = testData6[9544];
@(posedge clk);
#1;data_in = testData6[9545];
@(posedge clk);
#1;data_in = testData6[9546];
@(posedge clk);
#1;data_in = testData6[9547];
@(posedge clk);
#1;data_in = testData6[9548];
@(posedge clk);
#1;data_in = testData6[9549];
@(posedge clk);
#1;data_in = testData6[9550];
@(posedge clk);
#1;data_in = testData6[9551];
@(posedge clk);
#1;data_in = testData6[9552];
@(posedge clk);
#1;data_in = testData6[9553];
@(posedge clk);
#1;data_in = testData6[9554];
@(posedge clk);
#1;data_in = testData6[9555];
@(posedge clk);
#1;data_in = testData6[9556];
@(posedge clk);
#1;data_in = testData6[9557];
@(posedge clk);
#1;data_in = testData6[9558];
@(posedge clk);
#1;data_in = testData6[9559];
@(posedge clk);
#1;data_in = testData6[9560];
@(posedge clk);
#1;data_in = testData6[9561];
@(posedge clk);
#1;data_in = testData6[9562];
@(posedge clk);
#1;data_in = testData6[9563];
@(posedge clk);
#1;data_in = testData6[9564];
@(posedge clk);
#1;data_in = testData6[9565];
@(posedge clk);
#1;data_in = testData6[9566];
@(posedge clk);
#1;data_in = testData6[9567];
@(posedge clk);
#1;data_in = testData6[9568];
@(posedge clk);
#1;data_in = testData6[9569];
@(posedge clk);
#1;data_in = testData6[9570];
@(posedge clk);
#1;data_in = testData6[9571];
@(posedge clk);
#1;data_in = testData6[9572];
@(posedge clk);
#1;data_in = testData6[9573];
@(posedge clk);
#1;data_in = testData6[9574];
@(posedge clk);
#1;data_in = testData6[9575];
@(posedge clk);
#1;data_in = testData6[9576];
@(posedge clk);
#1;data_in = testData6[9577];
@(posedge clk);
#1;data_in = testData6[9578];
@(posedge clk);
#1;data_in = testData6[9579];
@(posedge clk);
#1;data_in = testData6[9580];
@(posedge clk);
#1;data_in = testData6[9581];
@(posedge clk);
#1;data_in = testData6[9582];
@(posedge clk);
#1;data_in = testData6[9583];
@(posedge clk);
#1;data_in = testData6[9584];
@(posedge clk);
#1;data_in = testData6[9585];
@(posedge clk);
#1;data_in = testData6[9586];
@(posedge clk);
#1;data_in = testData6[9587];
@(posedge clk);
#1;data_in = testData6[9588];
@(posedge clk);
#1;data_in = testData6[9589];
@(posedge clk);
#1;data_in = testData6[9590];
@(posedge clk);
#1;data_in = testData6[9591];
@(posedge clk);
#1;data_in = testData6[9592];
@(posedge clk);
#1;data_in = testData6[9593];
@(posedge clk);
#1;data_in = testData6[9594];
@(posedge clk);
#1;data_in = testData6[9595];
@(posedge clk);
#1;data_in = testData6[9596];
@(posedge clk);
#1;data_in = testData6[9597];
@(posedge clk);
#1;data_in = testData6[9598];
@(posedge clk);
#1;data_in = testData6[9599];
@(posedge clk);
#1;data_in = testData6[9600];
@(posedge clk);
#1;data_in = testData6[9601];
@(posedge clk);
#1;data_in = testData6[9602];
@(posedge clk);
#1;data_in = testData6[9603];
@(posedge clk);
#1;data_in = testData6[9604];
@(posedge clk);
#1;data_in = testData6[9605];
@(posedge clk);
#1;data_in = testData6[9606];
@(posedge clk);
#1;data_in = testData6[9607];
@(posedge clk);
#1;data_in = testData6[9608];
@(posedge clk);
#1;data_in = testData6[9609];
@(posedge clk);
#1;data_in = testData6[9610];
@(posedge clk);
#1;data_in = testData6[9611];
@(posedge clk);
#1;data_in = testData6[9612];
@(posedge clk);
#1;data_in = testData6[9613];
@(posedge clk);
#1;data_in = testData6[9614];
@(posedge clk);
#1;data_in = testData6[9615];
@(posedge clk);
#1;data_in = testData6[9616];
@(posedge clk);
#1;data_in = testData6[9617];
@(posedge clk);
#1;data_in = testData6[9618];
@(posedge clk);
#1;data_in = testData6[9619];
@(posedge clk);
#1;data_in = testData6[9620];
@(posedge clk);
#1;data_in = testData6[9621];
@(posedge clk);
#1;data_in = testData6[9622];
@(posedge clk);
#1;data_in = testData6[9623];
@(posedge clk);
#1;data_in = testData6[9624];
@(posedge clk);
#1;data_in = testData6[9625];
@(posedge clk);
#1;data_in = testData6[9626];
@(posedge clk);
#1;data_in = testData6[9627];
@(posedge clk);
#1;data_in = testData6[9628];
@(posedge clk);
#1;data_in = testData6[9629];
@(posedge clk);
#1;data_in = testData6[9630];
@(posedge clk);
#1;data_in = testData6[9631];
@(posedge clk);
#1;data_in = testData6[9632];
@(posedge clk);
#1;data_in = testData6[9633];
@(posedge clk);
#1;data_in = testData6[9634];
@(posedge clk);
#1;data_in = testData6[9635];
@(posedge clk);
#1;data_in = testData6[9636];
@(posedge clk);
#1;data_in = testData6[9637];
@(posedge clk);
#1;data_in = testData6[9638];
@(posedge clk);
#1;data_in = testData6[9639];
@(posedge clk);
#1;data_in = testData6[9640];
@(posedge clk);
#1;data_in = testData6[9641];
@(posedge clk);
#1;data_in = testData6[9642];
@(posedge clk);
#1;data_in = testData6[9643];
@(posedge clk);
#1;data_in = testData6[9644];
@(posedge clk);
#1;data_in = testData6[9645];
@(posedge clk);
#1;data_in = testData6[9646];
@(posedge clk);
#1;data_in = testData6[9647];
@(posedge clk);
#1;data_in = testData6[9648];
@(posedge clk);
#1;data_in = testData6[9649];
@(posedge clk);
#1;data_in = testData6[9650];
@(posedge clk);
#1;data_in = testData6[9651];
@(posedge clk);
#1;data_in = testData6[9652];
@(posedge clk);
#1;data_in = testData6[9653];
@(posedge clk);
#1;data_in = testData6[9654];
@(posedge clk);
#1;data_in = testData6[9655];
@(posedge clk);
#1;data_in = testData6[9656];
@(posedge clk);
#1;data_in = testData6[9657];
@(posedge clk);
#1;data_in = testData6[9658];
@(posedge clk);
#1;data_in = testData6[9659];
@(posedge clk);
#1;data_in = testData6[9660];
@(posedge clk);
#1;data_in = testData6[9661];
@(posedge clk);
#1;data_in = testData6[9662];
@(posedge clk);
#1;data_in = testData6[9663];
@(posedge clk);
#1;data_in = testData6[9664];
@(posedge clk);
#1;data_in = testData6[9665];
@(posedge clk);
#1;data_in = testData6[9666];
@(posedge clk);
#1;data_in = testData6[9667];
@(posedge clk);
#1;data_in = testData6[9668];
@(posedge clk);
#1;data_in = testData6[9669];
@(posedge clk);
#1;data_in = testData6[9670];
@(posedge clk);
#1;data_in = testData6[9671];
@(posedge clk);
#1;data_in = testData6[9672];
@(posedge clk);
#1;data_in = testData6[9673];
@(posedge clk);
#1;data_in = testData6[9674];
@(posedge clk);
#1;data_in = testData6[9675];
@(posedge clk);
#1;data_in = testData6[9676];
@(posedge clk);
#1;data_in = testData6[9677];
@(posedge clk);
#1;data_in = testData6[9678];
@(posedge clk);
#1;data_in = testData6[9679];
@(posedge clk);
#1;data_in = testData6[9680];
@(posedge clk);
#1;data_in = testData6[9681];
@(posedge clk);
#1;data_in = testData6[9682];
@(posedge clk);
#1;data_in = testData6[9683];
@(posedge clk);
#1;data_in = testData6[9684];
@(posedge clk);
#1;data_in = testData6[9685];
@(posedge clk);
#1;data_in = testData6[9686];
@(posedge clk);
#1;data_in = testData6[9687];
@(posedge clk);
#1;data_in = testData6[9688];
@(posedge clk);
#1;data_in = testData6[9689];
@(posedge clk);
#1;data_in = testData6[9690];
@(posedge clk);
#1;data_in = testData6[9691];
@(posedge clk);
#1;data_in = testData6[9692];
@(posedge clk);
#1;data_in = testData6[9693];
@(posedge clk);
#1;data_in = testData6[9694];
@(posedge clk);
#1;data_in = testData6[9695];
@(posedge clk);
#1;data_in = testData6[9696];
@(posedge clk);
#1;data_in = testData6[9697];
@(posedge clk);
#1;data_in = testData6[9698];
@(posedge clk);
#1;data_in = testData6[9699];
@(posedge clk);
#1;data_in = testData6[9700];
@(posedge clk);
#1;data_in = testData6[9701];
@(posedge clk);
#1;data_in = testData6[9702];
@(posedge clk);
#1;data_in = testData6[9703];
@(posedge clk);
#1;data_in = testData6[9704];
@(posedge clk);
#1;data_in = testData6[9705];
@(posedge clk);
#1;data_in = testData6[9706];
@(posedge clk);
#1;data_in = testData6[9707];
@(posedge clk);
#1;data_in = testData6[9708];
@(posedge clk);
#1;data_in = testData6[9709];
@(posedge clk);
#1;data_in = testData6[9710];
@(posedge clk);
#1;data_in = testData6[9711];
@(posedge clk);
#1;data_in = testData6[9712];
@(posedge clk);
#1;data_in = testData6[9713];
@(posedge clk);
#1;data_in = testData6[9714];
@(posedge clk);
#1;data_in = testData6[9715];
@(posedge clk);
#1;data_in = testData6[9716];
@(posedge clk);
#1;data_in = testData6[9717];
@(posedge clk);
#1;data_in = testData6[9718];
@(posedge clk);
#1;data_in = testData6[9719];
@(posedge clk);
#1;data_in = testData6[9720];
@(posedge clk);
#1;data_in = testData6[9721];
@(posedge clk);
#1;data_in = testData6[9722];
@(posedge clk);
#1;data_in = testData6[9723];
@(posedge clk);
#1;data_in = testData6[9724];
@(posedge clk);
#1;data_in = testData6[9725];
@(posedge clk);
#1;data_in = testData6[9726];
@(posedge clk);
#1;data_in = testData6[9727];
@(posedge clk);
#1;data_in = testData6[9728];
@(posedge clk);
#1;data_in = testData6[9729];
@(posedge clk);
#1;data_in = testData6[9730];
@(posedge clk);
#1;data_in = testData6[9731];
@(posedge clk);
#1;data_in = testData6[9732];
@(posedge clk);
#1;data_in = testData6[9733];
@(posedge clk);
#1;data_in = testData6[9734];
@(posedge clk);
#1;data_in = testData6[9735];
@(posedge clk);
#1;data_in = testData6[9736];
@(posedge clk);
#1;data_in = testData6[9737];
@(posedge clk);
#1;data_in = testData6[9738];
@(posedge clk);
#1;data_in = testData6[9739];
@(posedge clk);
#1;data_in = testData6[9740];
@(posedge clk);
#1;data_in = testData6[9741];
@(posedge clk);
#1;data_in = testData6[9742];
@(posedge clk);
#1;data_in = testData6[9743];
@(posedge clk);
#1;data_in = testData6[9744];
@(posedge clk);
#1;data_in = testData6[9745];
@(posedge clk);
#1;data_in = testData6[9746];
@(posedge clk);
#1;data_in = testData6[9747];
@(posedge clk);
#1;data_in = testData6[9748];
@(posedge clk);
#1;data_in = testData6[9749];
@(posedge clk);
#1;data_in = testData6[9750];
@(posedge clk);
#1;data_in = testData6[9751];
@(posedge clk);
#1;data_in = testData6[9752];
@(posedge clk);
#1;data_in = testData6[9753];
@(posedge clk);
#1;data_in = testData6[9754];
@(posedge clk);
#1;data_in = testData6[9755];
@(posedge clk);
#1;data_in = testData6[9756];
@(posedge clk);
#1;data_in = testData6[9757];
@(posedge clk);
#1;data_in = testData6[9758];
@(posedge clk);
#1;data_in = testData6[9759];
@(posedge clk);
#1;data_in = testData6[9760];
@(posedge clk);
#1;data_in = testData6[9761];
@(posedge clk);
#1;data_in = testData6[9762];
@(posedge clk);
#1;data_in = testData6[9763];
@(posedge clk);
#1;data_in = testData6[9764];
@(posedge clk);
#1;data_in = testData6[9765];
@(posedge clk);
#1;data_in = testData6[9766];
@(posedge clk);
#1;data_in = testData6[9767];
@(posedge clk);
#1;data_in = testData6[9768];
@(posedge clk);
#1;data_in = testData6[9769];
@(posedge clk);
#1;data_in = testData6[9770];
@(posedge clk);
#1;data_in = testData6[9771];
@(posedge clk);
#1;data_in = testData6[9772];
@(posedge clk);
#1;data_in = testData6[9773];
@(posedge clk);
#1;data_in = testData6[9774];
@(posedge clk);
#1;data_in = testData6[9775];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[9776]; 
@(posedge clk);
#1;data_in = testData6[9777];
@(posedge clk);
#1;data_in = testData6[9778];
@(posedge clk);
#1;data_in = testData6[9779];
@(posedge clk);
#1;data_in = testData6[9780];
@(posedge clk);
#1;data_in = testData6[9781];
@(posedge clk);
#1;data_in = testData6[9782];
@(posedge clk);
#1;data_in = testData6[9783];
@(posedge clk);
#1;data_in = testData6[9784];
@(posedge clk);
#1;data_in = testData6[9785];
@(posedge clk);
#1;data_in = testData6[9786];
@(posedge clk);
#1;data_in = testData6[9787];
@(posedge clk);
#1;data_in = testData6[9788];
@(posedge clk);
#1;data_in = testData6[9789];
@(posedge clk);
#1;data_in = testData6[9790];
@(posedge clk);
#1;data_in = testData6[9791];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[9792];
@(posedge clk);
#1;data_in = testData6[9793];
@(posedge clk);
#1;data_in = testData6[9794];
@(posedge clk);
#1;data_in = testData6[9795];
@(posedge clk);
#1;data_in = testData6[9796];
@(posedge clk);
#1;data_in = testData6[9797];
@(posedge clk);
#1;data_in = testData6[9798];
@(posedge clk);
#1;data_in = testData6[9799];
@(posedge clk);
#1;data_in = testData6[9800];
@(posedge clk);
#1;data_in = testData6[9801];
@(posedge clk);
#1;data_in = testData6[9802];
@(posedge clk);
#1;data_in = testData6[9803];
@(posedge clk);
#1;data_in = testData6[9804];
@(posedge clk);
#1;data_in = testData6[9805];
@(posedge clk);
#1;data_in = testData6[9806];
@(posedge clk);
#1;data_in = testData6[9807];
@(posedge clk);
#1;data_in = testData6[9808];
@(posedge clk);
#1;data_in = testData6[9809];
@(posedge clk);
#1;data_in = testData6[9810];
@(posedge clk);
#1;data_in = testData6[9811];
@(posedge clk);
#1;data_in = testData6[9812];
@(posedge clk);
#1;data_in = testData6[9813];
@(posedge clk);
#1;data_in = testData6[9814];
@(posedge clk);
#1;data_in = testData6[9815];
@(posedge clk);
#1;data_in = testData6[9816];
@(posedge clk);
#1;data_in = testData6[9817];
@(posedge clk);
#1;data_in = testData6[9818];
@(posedge clk);
#1;data_in = testData6[9819];
@(posedge clk);
#1;data_in = testData6[9820];
@(posedge clk);
#1;data_in = testData6[9821];
@(posedge clk);
#1;data_in = testData6[9822];
@(posedge clk);
#1;data_in = testData6[9823];
@(posedge clk);
#1;data_in = testData6[9824];
@(posedge clk);
#1;data_in = testData6[9825];
@(posedge clk);
#1;data_in = testData6[9826];
@(posedge clk);
#1;data_in = testData6[9827];
@(posedge clk);
#1;data_in = testData6[9828];
@(posedge clk);
#1;data_in = testData6[9829];
@(posedge clk);
#1;data_in = testData6[9830];
@(posedge clk);
#1;data_in = testData6[9831];
@(posedge clk);
#1;data_in = testData6[9832];
@(posedge clk);
#1;data_in = testData6[9833];
@(posedge clk);
#1;data_in = testData6[9834];
@(posedge clk);
#1;data_in = testData6[9835];
@(posedge clk);
#1;data_in = testData6[9836];
@(posedge clk);
#1;data_in = testData6[9837];
@(posedge clk);
#1;data_in = testData6[9838];
@(posedge clk);
#1;data_in = testData6[9839];
@(posedge clk);
#1;data_in = testData6[9840];
@(posedge clk);
#1;data_in = testData6[9841];
@(posedge clk);
#1;data_in = testData6[9842];
@(posedge clk);
#1;data_in = testData6[9843];
@(posedge clk);
#1;data_in = testData6[9844];
@(posedge clk);
#1;data_in = testData6[9845];
@(posedge clk);
#1;data_in = testData6[9846];
@(posedge clk);
#1;data_in = testData6[9847];
@(posedge clk);
#1;data_in = testData6[9848];
@(posedge clk);
#1;data_in = testData6[9849];
@(posedge clk);
#1;data_in = testData6[9850];
@(posedge clk);
#1;data_in = testData6[9851];
@(posedge clk);
#1;data_in = testData6[9852];
@(posedge clk);
#1;data_in = testData6[9853];
@(posedge clk);
#1;data_in = testData6[9854];
@(posedge clk);
#1;data_in = testData6[9855];
@(posedge clk);
#1;data_in = testData6[9856];
@(posedge clk);
#1;data_in = testData6[9857];
@(posedge clk);
#1;data_in = testData6[9858];
@(posedge clk);
#1;data_in = testData6[9859];
@(posedge clk);
#1;data_in = testData6[9860];
@(posedge clk);
#1;data_in = testData6[9861];
@(posedge clk);
#1;data_in = testData6[9862];
@(posedge clk);
#1;data_in = testData6[9863];
@(posedge clk);
#1;data_in = testData6[9864];
@(posedge clk);
#1;data_in = testData6[9865];
@(posedge clk);
#1;data_in = testData6[9866];
@(posedge clk);
#1;data_in = testData6[9867];
@(posedge clk);
#1;data_in = testData6[9868];
@(posedge clk);
#1;data_in = testData6[9869];
@(posedge clk);
#1;data_in = testData6[9870];
@(posedge clk);
#1;data_in = testData6[9871];
@(posedge clk);
#1;data_in = testData6[9872];
@(posedge clk);
#1;data_in = testData6[9873];
@(posedge clk);
#1;data_in = testData6[9874];
@(posedge clk);
#1;data_in = testData6[9875];
@(posedge clk);
#1;data_in = testData6[9876];
@(posedge clk);
#1;data_in = testData6[9877];
@(posedge clk);
#1;data_in = testData6[9878];
@(posedge clk);
#1;data_in = testData6[9879];
@(posedge clk);
#1;data_in = testData6[9880];
@(posedge clk);
#1;data_in = testData6[9881];
@(posedge clk);
#1;data_in = testData6[9882];
@(posedge clk);
#1;data_in = testData6[9883];
@(posedge clk);
#1;data_in = testData6[9884];
@(posedge clk);
#1;data_in = testData6[9885];
@(posedge clk);
#1;data_in = testData6[9886];
@(posedge clk);
#1;data_in = testData6[9887];
@(posedge clk);
#1;data_in = testData6[9888];
@(posedge clk);
#1;data_in = testData6[9889];
@(posedge clk);
#1;data_in = testData6[9890];
@(posedge clk);
#1;data_in = testData6[9891];
@(posedge clk);
#1;data_in = testData6[9892];
@(posedge clk);
#1;data_in = testData6[9893];
@(posedge clk);
#1;data_in = testData6[9894];
@(posedge clk);
#1;data_in = testData6[9895];
@(posedge clk);
#1;data_in = testData6[9896];
@(posedge clk);
#1;data_in = testData6[9897];
@(posedge clk);
#1;data_in = testData6[9898];
@(posedge clk);
#1;data_in = testData6[9899];
@(posedge clk);
#1;data_in = testData6[9900];
@(posedge clk);
#1;data_in = testData6[9901];
@(posedge clk);
#1;data_in = testData6[9902];
@(posedge clk);
#1;data_in = testData6[9903];
@(posedge clk);
#1;data_in = testData6[9904];
@(posedge clk);
#1;data_in = testData6[9905];
@(posedge clk);
#1;data_in = testData6[9906];
@(posedge clk);
#1;data_in = testData6[9907];
@(posedge clk);
#1;data_in = testData6[9908];
@(posedge clk);
#1;data_in = testData6[9909];
@(posedge clk);
#1;data_in = testData6[9910];
@(posedge clk);
#1;data_in = testData6[9911];
@(posedge clk);
#1;data_in = testData6[9912];
@(posedge clk);
#1;data_in = testData6[9913];
@(posedge clk);
#1;data_in = testData6[9914];
@(posedge clk);
#1;data_in = testData6[9915];
@(posedge clk);
#1;data_in = testData6[9916];
@(posedge clk);
#1;data_in = testData6[9917];
@(posedge clk);
#1;data_in = testData6[9918];
@(posedge clk);
#1;data_in = testData6[9919];
@(posedge clk);
#1;data_in = testData6[9920];
@(posedge clk);
#1;data_in = testData6[9921];
@(posedge clk);
#1;data_in = testData6[9922];
@(posedge clk);
#1;data_in = testData6[9923];
@(posedge clk);
#1;data_in = testData6[9924];
@(posedge clk);
#1;data_in = testData6[9925];
@(posedge clk);
#1;data_in = testData6[9926];
@(posedge clk);
#1;data_in = testData6[9927];
@(posedge clk);
#1;data_in = testData6[9928];
@(posedge clk);
#1;data_in = testData6[9929];
@(posedge clk);
#1;data_in = testData6[9930];
@(posedge clk);
#1;data_in = testData6[9931];
@(posedge clk);
#1;data_in = testData6[9932];
@(posedge clk);
#1;data_in = testData6[9933];
@(posedge clk);
#1;data_in = testData6[9934];
@(posedge clk);
#1;data_in = testData6[9935];
@(posedge clk);
#1;data_in = testData6[9936];
@(posedge clk);
#1;data_in = testData6[9937];
@(posedge clk);
#1;data_in = testData6[9938];
@(posedge clk);
#1;data_in = testData6[9939];
@(posedge clk);
#1;data_in = testData6[9940];
@(posedge clk);
#1;data_in = testData6[9941];
@(posedge clk);
#1;data_in = testData6[9942];
@(posedge clk);
#1;data_in = testData6[9943];
@(posedge clk);
#1;data_in = testData6[9944];
@(posedge clk);
#1;data_in = testData6[9945];
@(posedge clk);
#1;data_in = testData6[9946];
@(posedge clk);
#1;data_in = testData6[9947];
@(posedge clk);
#1;data_in = testData6[9948];
@(posedge clk);
#1;data_in = testData6[9949];
@(posedge clk);
#1;data_in = testData6[9950];
@(posedge clk);
#1;data_in = testData6[9951];
@(posedge clk);
#1;data_in = testData6[9952];
@(posedge clk);
#1;data_in = testData6[9953];
@(posedge clk);
#1;data_in = testData6[9954];
@(posedge clk);
#1;data_in = testData6[9955];
@(posedge clk);
#1;data_in = testData6[9956];
@(posedge clk);
#1;data_in = testData6[9957];
@(posedge clk);
#1;data_in = testData6[9958];
@(posedge clk);
#1;data_in = testData6[9959];
@(posedge clk);
#1;data_in = testData6[9960];
@(posedge clk);
#1;data_in = testData6[9961];
@(posedge clk);
#1;data_in = testData6[9962];
@(posedge clk);
#1;data_in = testData6[9963];
@(posedge clk);
#1;data_in = testData6[9964];
@(posedge clk);
#1;data_in = testData6[9965];
@(posedge clk);
#1;data_in = testData6[9966];
@(posedge clk);
#1;data_in = testData6[9967];
@(posedge clk);
#1;data_in = testData6[9968];
@(posedge clk);
#1;data_in = testData6[9969];
@(posedge clk);
#1;data_in = testData6[9970];
@(posedge clk);
#1;data_in = testData6[9971];
@(posedge clk);
#1;data_in = testData6[9972];
@(posedge clk);
#1;data_in = testData6[9973];
@(posedge clk);
#1;data_in = testData6[9974];
@(posedge clk);
#1;data_in = testData6[9975];
@(posedge clk);
#1;data_in = testData6[9976];
@(posedge clk);
#1;data_in = testData6[9977];
@(posedge clk);
#1;data_in = testData6[9978];
@(posedge clk);
#1;data_in = testData6[9979];
@(posedge clk);
#1;data_in = testData6[9980];
@(posedge clk);
#1;data_in = testData6[9981];
@(posedge clk);
#1;data_in = testData6[9982];
@(posedge clk);
#1;data_in = testData6[9983];
@(posedge clk);
#1;data_in = testData6[9984];
@(posedge clk);
#1;data_in = testData6[9985];
@(posedge clk);
#1;data_in = testData6[9986];
@(posedge clk);
#1;data_in = testData6[9987];
@(posedge clk);
#1;data_in = testData6[9988];
@(posedge clk);
#1;data_in = testData6[9989];
@(posedge clk);
#1;data_in = testData6[9990];
@(posedge clk);
#1;data_in = testData6[9991];
@(posedge clk);
#1;data_in = testData6[9992];
@(posedge clk);
#1;data_in = testData6[9993];
@(posedge clk);
#1;data_in = testData6[9994];
@(posedge clk);
#1;data_in = testData6[9995];
@(posedge clk);
#1;data_in = testData6[9996];
@(posedge clk);
#1;data_in = testData6[9997];
@(posedge clk);
#1;data_in = testData6[9998];
@(posedge clk);
#1;data_in = testData6[9999];
@(posedge clk);
#1;data_in = testData6[10000];
@(posedge clk);
#1;data_in = testData6[10001];
@(posedge clk);
#1;data_in = testData6[10002];
@(posedge clk);
#1;data_in = testData6[10003];
@(posedge clk);
#1;data_in = testData6[10004];
@(posedge clk);
#1;data_in = testData6[10005];
@(posedge clk);
#1;data_in = testData6[10006];
@(posedge clk);
#1;data_in = testData6[10007];
@(posedge clk);
#1;data_in = testData6[10008];
@(posedge clk);
#1;data_in = testData6[10009];
@(posedge clk);
#1;data_in = testData6[10010];
@(posedge clk);
#1;data_in = testData6[10011];
@(posedge clk);
#1;data_in = testData6[10012];
@(posedge clk);
#1;data_in = testData6[10013];
@(posedge clk);
#1;data_in = testData6[10014];
@(posedge clk);
#1;data_in = testData6[10015];
@(posedge clk);
#1;data_in = testData6[10016];
@(posedge clk);
#1;data_in = testData6[10017];
@(posedge clk);
#1;data_in = testData6[10018];
@(posedge clk);
#1;data_in = testData6[10019];
@(posedge clk);
#1;data_in = testData6[10020];
@(posedge clk);
#1;data_in = testData6[10021];
@(posedge clk);
#1;data_in = testData6[10022];
@(posedge clk);
#1;data_in = testData6[10023];
@(posedge clk);
#1;data_in = testData6[10024];
@(posedge clk);
#1;data_in = testData6[10025];
@(posedge clk);
#1;data_in = testData6[10026];
@(posedge clk);
#1;data_in = testData6[10027];
@(posedge clk);
#1;data_in = testData6[10028];
@(posedge clk);
#1;data_in = testData6[10029];
@(posedge clk);
#1;data_in = testData6[10030];
@(posedge clk);
#1;data_in = testData6[10031];
@(posedge clk);
#1;data_in = testData6[10032];
@(posedge clk);
#1;data_in = testData6[10033];
@(posedge clk);
#1;data_in = testData6[10034];
@(posedge clk);
#1;data_in = testData6[10035];
@(posedge clk);
#1;data_in = testData6[10036];
@(posedge clk);
#1;data_in = testData6[10037];
@(posedge clk);
#1;data_in = testData6[10038];
@(posedge clk);
#1;data_in = testData6[10039];
@(posedge clk);
#1;data_in = testData6[10040];
@(posedge clk);
#1;data_in = testData6[10041];
@(posedge clk);
#1;data_in = testData6[10042];
@(posedge clk);
#1;data_in = testData6[10043];
@(posedge clk);
#1;data_in = testData6[10044];
@(posedge clk);
#1;data_in = testData6[10045];
@(posedge clk);
#1;data_in = testData6[10046];
@(posedge clk);
#1;data_in = testData6[10047];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[10048]; 
@(posedge clk);
#1;data_in = testData6[10049];
@(posedge clk);
#1;data_in = testData6[10050];
@(posedge clk);
#1;data_in = testData6[10051];
@(posedge clk);
#1;data_in = testData6[10052];
@(posedge clk);
#1;data_in = testData6[10053];
@(posedge clk);
#1;data_in = testData6[10054];
@(posedge clk);
#1;data_in = testData6[10055];
@(posedge clk);
#1;data_in = testData6[10056];
@(posedge clk);
#1;data_in = testData6[10057];
@(posedge clk);
#1;data_in = testData6[10058];
@(posedge clk);
#1;data_in = testData6[10059];
@(posedge clk);
#1;data_in = testData6[10060];
@(posedge clk);
#1;data_in = testData6[10061];
@(posedge clk);
#1;data_in = testData6[10062];
@(posedge clk);
#1;data_in = testData6[10063];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[10064];
@(posedge clk);
#1;data_in = testData6[10065];
@(posedge clk);
#1;data_in = testData6[10066];
@(posedge clk);
#1;data_in = testData6[10067];
@(posedge clk);
#1;data_in = testData6[10068];
@(posedge clk);
#1;data_in = testData6[10069];
@(posedge clk);
#1;data_in = testData6[10070];
@(posedge clk);
#1;data_in = testData6[10071];
@(posedge clk);
#1;data_in = testData6[10072];
@(posedge clk);
#1;data_in = testData6[10073];
@(posedge clk);
#1;data_in = testData6[10074];
@(posedge clk);
#1;data_in = testData6[10075];
@(posedge clk);
#1;data_in = testData6[10076];
@(posedge clk);
#1;data_in = testData6[10077];
@(posedge clk);
#1;data_in = testData6[10078];
@(posedge clk);
#1;data_in = testData6[10079];
@(posedge clk);
#1;data_in = testData6[10080];
@(posedge clk);
#1;data_in = testData6[10081];
@(posedge clk);
#1;data_in = testData6[10082];
@(posedge clk);
#1;data_in = testData6[10083];
@(posedge clk);
#1;data_in = testData6[10084];
@(posedge clk);
#1;data_in = testData6[10085];
@(posedge clk);
#1;data_in = testData6[10086];
@(posedge clk);
#1;data_in = testData6[10087];
@(posedge clk);
#1;data_in = testData6[10088];
@(posedge clk);
#1;data_in = testData6[10089];
@(posedge clk);
#1;data_in = testData6[10090];
@(posedge clk);
#1;data_in = testData6[10091];
@(posedge clk);
#1;data_in = testData6[10092];
@(posedge clk);
#1;data_in = testData6[10093];
@(posedge clk);
#1;data_in = testData6[10094];
@(posedge clk);
#1;data_in = testData6[10095];
@(posedge clk);
#1;data_in = testData6[10096];
@(posedge clk);
#1;data_in = testData6[10097];
@(posedge clk);
#1;data_in = testData6[10098];
@(posedge clk);
#1;data_in = testData6[10099];
@(posedge clk);
#1;data_in = testData6[10100];
@(posedge clk);
#1;data_in = testData6[10101];
@(posedge clk);
#1;data_in = testData6[10102];
@(posedge clk);
#1;data_in = testData6[10103];
@(posedge clk);
#1;data_in = testData6[10104];
@(posedge clk);
#1;data_in = testData6[10105];
@(posedge clk);
#1;data_in = testData6[10106];
@(posedge clk);
#1;data_in = testData6[10107];
@(posedge clk);
#1;data_in = testData6[10108];
@(posedge clk);
#1;data_in = testData6[10109];
@(posedge clk);
#1;data_in = testData6[10110];
@(posedge clk);
#1;data_in = testData6[10111];
@(posedge clk);
#1;data_in = testData6[10112];
@(posedge clk);
#1;data_in = testData6[10113];
@(posedge clk);
#1;data_in = testData6[10114];
@(posedge clk);
#1;data_in = testData6[10115];
@(posedge clk);
#1;data_in = testData6[10116];
@(posedge clk);
#1;data_in = testData6[10117];
@(posedge clk);
#1;data_in = testData6[10118];
@(posedge clk);
#1;data_in = testData6[10119];
@(posedge clk);
#1;data_in = testData6[10120];
@(posedge clk);
#1;data_in = testData6[10121];
@(posedge clk);
#1;data_in = testData6[10122];
@(posedge clk);
#1;data_in = testData6[10123];
@(posedge clk);
#1;data_in = testData6[10124];
@(posedge clk);
#1;data_in = testData6[10125];
@(posedge clk);
#1;data_in = testData6[10126];
@(posedge clk);
#1;data_in = testData6[10127];
@(posedge clk);
#1;data_in = testData6[10128];
@(posedge clk);
#1;data_in = testData6[10129];
@(posedge clk);
#1;data_in = testData6[10130];
@(posedge clk);
#1;data_in = testData6[10131];
@(posedge clk);
#1;data_in = testData6[10132];
@(posedge clk);
#1;data_in = testData6[10133];
@(posedge clk);
#1;data_in = testData6[10134];
@(posedge clk);
#1;data_in = testData6[10135];
@(posedge clk);
#1;data_in = testData6[10136];
@(posedge clk);
#1;data_in = testData6[10137];
@(posedge clk);
#1;data_in = testData6[10138];
@(posedge clk);
#1;data_in = testData6[10139];
@(posedge clk);
#1;data_in = testData6[10140];
@(posedge clk);
#1;data_in = testData6[10141];
@(posedge clk);
#1;data_in = testData6[10142];
@(posedge clk);
#1;data_in = testData6[10143];
@(posedge clk);
#1;data_in = testData6[10144];
@(posedge clk);
#1;data_in = testData6[10145];
@(posedge clk);
#1;data_in = testData6[10146];
@(posedge clk);
#1;data_in = testData6[10147];
@(posedge clk);
#1;data_in = testData6[10148];
@(posedge clk);
#1;data_in = testData6[10149];
@(posedge clk);
#1;data_in = testData6[10150];
@(posedge clk);
#1;data_in = testData6[10151];
@(posedge clk);
#1;data_in = testData6[10152];
@(posedge clk);
#1;data_in = testData6[10153];
@(posedge clk);
#1;data_in = testData6[10154];
@(posedge clk);
#1;data_in = testData6[10155];
@(posedge clk);
#1;data_in = testData6[10156];
@(posedge clk);
#1;data_in = testData6[10157];
@(posedge clk);
#1;data_in = testData6[10158];
@(posedge clk);
#1;data_in = testData6[10159];
@(posedge clk);
#1;data_in = testData6[10160];
@(posedge clk);
#1;data_in = testData6[10161];
@(posedge clk);
#1;data_in = testData6[10162];
@(posedge clk);
#1;data_in = testData6[10163];
@(posedge clk);
#1;data_in = testData6[10164];
@(posedge clk);
#1;data_in = testData6[10165];
@(posedge clk);
#1;data_in = testData6[10166];
@(posedge clk);
#1;data_in = testData6[10167];
@(posedge clk);
#1;data_in = testData6[10168];
@(posedge clk);
#1;data_in = testData6[10169];
@(posedge clk);
#1;data_in = testData6[10170];
@(posedge clk);
#1;data_in = testData6[10171];
@(posedge clk);
#1;data_in = testData6[10172];
@(posedge clk);
#1;data_in = testData6[10173];
@(posedge clk);
#1;data_in = testData6[10174];
@(posedge clk);
#1;data_in = testData6[10175];
@(posedge clk);
#1;data_in = testData6[10176];
@(posedge clk);
#1;data_in = testData6[10177];
@(posedge clk);
#1;data_in = testData6[10178];
@(posedge clk);
#1;data_in = testData6[10179];
@(posedge clk);
#1;data_in = testData6[10180];
@(posedge clk);
#1;data_in = testData6[10181];
@(posedge clk);
#1;data_in = testData6[10182];
@(posedge clk);
#1;data_in = testData6[10183];
@(posedge clk);
#1;data_in = testData6[10184];
@(posedge clk);
#1;data_in = testData6[10185];
@(posedge clk);
#1;data_in = testData6[10186];
@(posedge clk);
#1;data_in = testData6[10187];
@(posedge clk);
#1;data_in = testData6[10188];
@(posedge clk);
#1;data_in = testData6[10189];
@(posedge clk);
#1;data_in = testData6[10190];
@(posedge clk);
#1;data_in = testData6[10191];
@(posedge clk);
#1;data_in = testData6[10192];
@(posedge clk);
#1;data_in = testData6[10193];
@(posedge clk);
#1;data_in = testData6[10194];
@(posedge clk);
#1;data_in = testData6[10195];
@(posedge clk);
#1;data_in = testData6[10196];
@(posedge clk);
#1;data_in = testData6[10197];
@(posedge clk);
#1;data_in = testData6[10198];
@(posedge clk);
#1;data_in = testData6[10199];
@(posedge clk);
#1;data_in = testData6[10200];
@(posedge clk);
#1;data_in = testData6[10201];
@(posedge clk);
#1;data_in = testData6[10202];
@(posedge clk);
#1;data_in = testData6[10203];
@(posedge clk);
#1;data_in = testData6[10204];
@(posedge clk);
#1;data_in = testData6[10205];
@(posedge clk);
#1;data_in = testData6[10206];
@(posedge clk);
#1;data_in = testData6[10207];
@(posedge clk);
#1;data_in = testData6[10208];
@(posedge clk);
#1;data_in = testData6[10209];
@(posedge clk);
#1;data_in = testData6[10210];
@(posedge clk);
#1;data_in = testData6[10211];
@(posedge clk);
#1;data_in = testData6[10212];
@(posedge clk);
#1;data_in = testData6[10213];
@(posedge clk);
#1;data_in = testData6[10214];
@(posedge clk);
#1;data_in = testData6[10215];
@(posedge clk);
#1;data_in = testData6[10216];
@(posedge clk);
#1;data_in = testData6[10217];
@(posedge clk);
#1;data_in = testData6[10218];
@(posedge clk);
#1;data_in = testData6[10219];
@(posedge clk);
#1;data_in = testData6[10220];
@(posedge clk);
#1;data_in = testData6[10221];
@(posedge clk);
#1;data_in = testData6[10222];
@(posedge clk);
#1;data_in = testData6[10223];
@(posedge clk);
#1;data_in = testData6[10224];
@(posedge clk);
#1;data_in = testData6[10225];
@(posedge clk);
#1;data_in = testData6[10226];
@(posedge clk);
#1;data_in = testData6[10227];
@(posedge clk);
#1;data_in = testData6[10228];
@(posedge clk);
#1;data_in = testData6[10229];
@(posedge clk);
#1;data_in = testData6[10230];
@(posedge clk);
#1;data_in = testData6[10231];
@(posedge clk);
#1;data_in = testData6[10232];
@(posedge clk);
#1;data_in = testData6[10233];
@(posedge clk);
#1;data_in = testData6[10234];
@(posedge clk);
#1;data_in = testData6[10235];
@(posedge clk);
#1;data_in = testData6[10236];
@(posedge clk);
#1;data_in = testData6[10237];
@(posedge clk);
#1;data_in = testData6[10238];
@(posedge clk);
#1;data_in = testData6[10239];
@(posedge clk);
#1;data_in = testData6[10240];
@(posedge clk);
#1;data_in = testData6[10241];
@(posedge clk);
#1;data_in = testData6[10242];
@(posedge clk);
#1;data_in = testData6[10243];
@(posedge clk);
#1;data_in = testData6[10244];
@(posedge clk);
#1;data_in = testData6[10245];
@(posedge clk);
#1;data_in = testData6[10246];
@(posedge clk);
#1;data_in = testData6[10247];
@(posedge clk);
#1;data_in = testData6[10248];
@(posedge clk);
#1;data_in = testData6[10249];
@(posedge clk);
#1;data_in = testData6[10250];
@(posedge clk);
#1;data_in = testData6[10251];
@(posedge clk);
#1;data_in = testData6[10252];
@(posedge clk);
#1;data_in = testData6[10253];
@(posedge clk);
#1;data_in = testData6[10254];
@(posedge clk);
#1;data_in = testData6[10255];
@(posedge clk);
#1;data_in = testData6[10256];
@(posedge clk);
#1;data_in = testData6[10257];
@(posedge clk);
#1;data_in = testData6[10258];
@(posedge clk);
#1;data_in = testData6[10259];
@(posedge clk);
#1;data_in = testData6[10260];
@(posedge clk);
#1;data_in = testData6[10261];
@(posedge clk);
#1;data_in = testData6[10262];
@(posedge clk);
#1;data_in = testData6[10263];
@(posedge clk);
#1;data_in = testData6[10264];
@(posedge clk);
#1;data_in = testData6[10265];
@(posedge clk);
#1;data_in = testData6[10266];
@(posedge clk);
#1;data_in = testData6[10267];
@(posedge clk);
#1;data_in = testData6[10268];
@(posedge clk);
#1;data_in = testData6[10269];
@(posedge clk);
#1;data_in = testData6[10270];
@(posedge clk);
#1;data_in = testData6[10271];
@(posedge clk);
#1;data_in = testData6[10272];
@(posedge clk);
#1;data_in = testData6[10273];
@(posedge clk);
#1;data_in = testData6[10274];
@(posedge clk);
#1;data_in = testData6[10275];
@(posedge clk);
#1;data_in = testData6[10276];
@(posedge clk);
#1;data_in = testData6[10277];
@(posedge clk);
#1;data_in = testData6[10278];
@(posedge clk);
#1;data_in = testData6[10279];
@(posedge clk);
#1;data_in = testData6[10280];
@(posedge clk);
#1;data_in = testData6[10281];
@(posedge clk);
#1;data_in = testData6[10282];
@(posedge clk);
#1;data_in = testData6[10283];
@(posedge clk);
#1;data_in = testData6[10284];
@(posedge clk);
#1;data_in = testData6[10285];
@(posedge clk);
#1;data_in = testData6[10286];
@(posedge clk);
#1;data_in = testData6[10287];
@(posedge clk);
#1;data_in = testData6[10288];
@(posedge clk);
#1;data_in = testData6[10289];
@(posedge clk);
#1;data_in = testData6[10290];
@(posedge clk);
#1;data_in = testData6[10291];
@(posedge clk);
#1;data_in = testData6[10292];
@(posedge clk);
#1;data_in = testData6[10293];
@(posedge clk);
#1;data_in = testData6[10294];
@(posedge clk);
#1;data_in = testData6[10295];
@(posedge clk);
#1;data_in = testData6[10296];
@(posedge clk);
#1;data_in = testData6[10297];
@(posedge clk);
#1;data_in = testData6[10298];
@(posedge clk);
#1;data_in = testData6[10299];
@(posedge clk);
#1;data_in = testData6[10300];
@(posedge clk);
#1;data_in = testData6[10301];
@(posedge clk);
#1;data_in = testData6[10302];
@(posedge clk);
#1;data_in = testData6[10303];
@(posedge clk);
#1;data_in = testData6[10304];
@(posedge clk);
#1;data_in = testData6[10305];
@(posedge clk);
#1;data_in = testData6[10306];
@(posedge clk);
#1;data_in = testData6[10307];
@(posedge clk);
#1;data_in = testData6[10308];
@(posedge clk);
#1;data_in = testData6[10309];
@(posedge clk);
#1;data_in = testData6[10310];
@(posedge clk);
#1;data_in = testData6[10311];
@(posedge clk);
#1;data_in = testData6[10312];
@(posedge clk);
#1;data_in = testData6[10313];
@(posedge clk);
#1;data_in = testData6[10314];
@(posedge clk);
#1;data_in = testData6[10315];
@(posedge clk);
#1;data_in = testData6[10316];
@(posedge clk);
#1;data_in = testData6[10317];
@(posedge clk);
#1;data_in = testData6[10318];
@(posedge clk);
#1;data_in = testData6[10319];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[10320]; 
@(posedge clk);
#1;data_in = testData6[10321];
@(posedge clk);
#1;data_in = testData6[10322];
@(posedge clk);
#1;data_in = testData6[10323];
@(posedge clk);
#1;data_in = testData6[10324];
@(posedge clk);
#1;data_in = testData6[10325];
@(posedge clk);
#1;data_in = testData6[10326];
@(posedge clk);
#1;data_in = testData6[10327];
@(posedge clk);
#1;data_in = testData6[10328];
@(posedge clk);
#1;data_in = testData6[10329];
@(posedge clk);
#1;data_in = testData6[10330];
@(posedge clk);
#1;data_in = testData6[10331];
@(posedge clk);
#1;data_in = testData6[10332];
@(posedge clk);
#1;data_in = testData6[10333];
@(posedge clk);
#1;data_in = testData6[10334];
@(posedge clk);
#1;data_in = testData6[10335];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[10336];
@(posedge clk);
#1;data_in = testData6[10337];
@(posedge clk);
#1;data_in = testData6[10338];
@(posedge clk);
#1;data_in = testData6[10339];
@(posedge clk);
#1;data_in = testData6[10340];
@(posedge clk);
#1;data_in = testData6[10341];
@(posedge clk);
#1;data_in = testData6[10342];
@(posedge clk);
#1;data_in = testData6[10343];
@(posedge clk);
#1;data_in = testData6[10344];
@(posedge clk);
#1;data_in = testData6[10345];
@(posedge clk);
#1;data_in = testData6[10346];
@(posedge clk);
#1;data_in = testData6[10347];
@(posedge clk);
#1;data_in = testData6[10348];
@(posedge clk);
#1;data_in = testData6[10349];
@(posedge clk);
#1;data_in = testData6[10350];
@(posedge clk);
#1;data_in = testData6[10351];
@(posedge clk);
#1;data_in = testData6[10352];
@(posedge clk);
#1;data_in = testData6[10353];
@(posedge clk);
#1;data_in = testData6[10354];
@(posedge clk);
#1;data_in = testData6[10355];
@(posedge clk);
#1;data_in = testData6[10356];
@(posedge clk);
#1;data_in = testData6[10357];
@(posedge clk);
#1;data_in = testData6[10358];
@(posedge clk);
#1;data_in = testData6[10359];
@(posedge clk);
#1;data_in = testData6[10360];
@(posedge clk);
#1;data_in = testData6[10361];
@(posedge clk);
#1;data_in = testData6[10362];
@(posedge clk);
#1;data_in = testData6[10363];
@(posedge clk);
#1;data_in = testData6[10364];
@(posedge clk);
#1;data_in = testData6[10365];
@(posedge clk);
#1;data_in = testData6[10366];
@(posedge clk);
#1;data_in = testData6[10367];
@(posedge clk);
#1;data_in = testData6[10368];
@(posedge clk);
#1;data_in = testData6[10369];
@(posedge clk);
#1;data_in = testData6[10370];
@(posedge clk);
#1;data_in = testData6[10371];
@(posedge clk);
#1;data_in = testData6[10372];
@(posedge clk);
#1;data_in = testData6[10373];
@(posedge clk);
#1;data_in = testData6[10374];
@(posedge clk);
#1;data_in = testData6[10375];
@(posedge clk);
#1;data_in = testData6[10376];
@(posedge clk);
#1;data_in = testData6[10377];
@(posedge clk);
#1;data_in = testData6[10378];
@(posedge clk);
#1;data_in = testData6[10379];
@(posedge clk);
#1;data_in = testData6[10380];
@(posedge clk);
#1;data_in = testData6[10381];
@(posedge clk);
#1;data_in = testData6[10382];
@(posedge clk);
#1;data_in = testData6[10383];
@(posedge clk);
#1;data_in = testData6[10384];
@(posedge clk);
#1;data_in = testData6[10385];
@(posedge clk);
#1;data_in = testData6[10386];
@(posedge clk);
#1;data_in = testData6[10387];
@(posedge clk);
#1;data_in = testData6[10388];
@(posedge clk);
#1;data_in = testData6[10389];
@(posedge clk);
#1;data_in = testData6[10390];
@(posedge clk);
#1;data_in = testData6[10391];
@(posedge clk);
#1;data_in = testData6[10392];
@(posedge clk);
#1;data_in = testData6[10393];
@(posedge clk);
#1;data_in = testData6[10394];
@(posedge clk);
#1;data_in = testData6[10395];
@(posedge clk);
#1;data_in = testData6[10396];
@(posedge clk);
#1;data_in = testData6[10397];
@(posedge clk);
#1;data_in = testData6[10398];
@(posedge clk);
#1;data_in = testData6[10399];
@(posedge clk);
#1;data_in = testData6[10400];
@(posedge clk);
#1;data_in = testData6[10401];
@(posedge clk);
#1;data_in = testData6[10402];
@(posedge clk);
#1;data_in = testData6[10403];
@(posedge clk);
#1;data_in = testData6[10404];
@(posedge clk);
#1;data_in = testData6[10405];
@(posedge clk);
#1;data_in = testData6[10406];
@(posedge clk);
#1;data_in = testData6[10407];
@(posedge clk);
#1;data_in = testData6[10408];
@(posedge clk);
#1;data_in = testData6[10409];
@(posedge clk);
#1;data_in = testData6[10410];
@(posedge clk);
#1;data_in = testData6[10411];
@(posedge clk);
#1;data_in = testData6[10412];
@(posedge clk);
#1;data_in = testData6[10413];
@(posedge clk);
#1;data_in = testData6[10414];
@(posedge clk);
#1;data_in = testData6[10415];
@(posedge clk);
#1;data_in = testData6[10416];
@(posedge clk);
#1;data_in = testData6[10417];
@(posedge clk);
#1;data_in = testData6[10418];
@(posedge clk);
#1;data_in = testData6[10419];
@(posedge clk);
#1;data_in = testData6[10420];
@(posedge clk);
#1;data_in = testData6[10421];
@(posedge clk);
#1;data_in = testData6[10422];
@(posedge clk);
#1;data_in = testData6[10423];
@(posedge clk);
#1;data_in = testData6[10424];
@(posedge clk);
#1;data_in = testData6[10425];
@(posedge clk);
#1;data_in = testData6[10426];
@(posedge clk);
#1;data_in = testData6[10427];
@(posedge clk);
#1;data_in = testData6[10428];
@(posedge clk);
#1;data_in = testData6[10429];
@(posedge clk);
#1;data_in = testData6[10430];
@(posedge clk);
#1;data_in = testData6[10431];
@(posedge clk);
#1;data_in = testData6[10432];
@(posedge clk);
#1;data_in = testData6[10433];
@(posedge clk);
#1;data_in = testData6[10434];
@(posedge clk);
#1;data_in = testData6[10435];
@(posedge clk);
#1;data_in = testData6[10436];
@(posedge clk);
#1;data_in = testData6[10437];
@(posedge clk);
#1;data_in = testData6[10438];
@(posedge clk);
#1;data_in = testData6[10439];
@(posedge clk);
#1;data_in = testData6[10440];
@(posedge clk);
#1;data_in = testData6[10441];
@(posedge clk);
#1;data_in = testData6[10442];
@(posedge clk);
#1;data_in = testData6[10443];
@(posedge clk);
#1;data_in = testData6[10444];
@(posedge clk);
#1;data_in = testData6[10445];
@(posedge clk);
#1;data_in = testData6[10446];
@(posedge clk);
#1;data_in = testData6[10447];
@(posedge clk);
#1;data_in = testData6[10448];
@(posedge clk);
#1;data_in = testData6[10449];
@(posedge clk);
#1;data_in = testData6[10450];
@(posedge clk);
#1;data_in = testData6[10451];
@(posedge clk);
#1;data_in = testData6[10452];
@(posedge clk);
#1;data_in = testData6[10453];
@(posedge clk);
#1;data_in = testData6[10454];
@(posedge clk);
#1;data_in = testData6[10455];
@(posedge clk);
#1;data_in = testData6[10456];
@(posedge clk);
#1;data_in = testData6[10457];
@(posedge clk);
#1;data_in = testData6[10458];
@(posedge clk);
#1;data_in = testData6[10459];
@(posedge clk);
#1;data_in = testData6[10460];
@(posedge clk);
#1;data_in = testData6[10461];
@(posedge clk);
#1;data_in = testData6[10462];
@(posedge clk);
#1;data_in = testData6[10463];
@(posedge clk);
#1;data_in = testData6[10464];
@(posedge clk);
#1;data_in = testData6[10465];
@(posedge clk);
#1;data_in = testData6[10466];
@(posedge clk);
#1;data_in = testData6[10467];
@(posedge clk);
#1;data_in = testData6[10468];
@(posedge clk);
#1;data_in = testData6[10469];
@(posedge clk);
#1;data_in = testData6[10470];
@(posedge clk);
#1;data_in = testData6[10471];
@(posedge clk);
#1;data_in = testData6[10472];
@(posedge clk);
#1;data_in = testData6[10473];
@(posedge clk);
#1;data_in = testData6[10474];
@(posedge clk);
#1;data_in = testData6[10475];
@(posedge clk);
#1;data_in = testData6[10476];
@(posedge clk);
#1;data_in = testData6[10477];
@(posedge clk);
#1;data_in = testData6[10478];
@(posedge clk);
#1;data_in = testData6[10479];
@(posedge clk);
#1;data_in = testData6[10480];
@(posedge clk);
#1;data_in = testData6[10481];
@(posedge clk);
#1;data_in = testData6[10482];
@(posedge clk);
#1;data_in = testData6[10483];
@(posedge clk);
#1;data_in = testData6[10484];
@(posedge clk);
#1;data_in = testData6[10485];
@(posedge clk);
#1;data_in = testData6[10486];
@(posedge clk);
#1;data_in = testData6[10487];
@(posedge clk);
#1;data_in = testData6[10488];
@(posedge clk);
#1;data_in = testData6[10489];
@(posedge clk);
#1;data_in = testData6[10490];
@(posedge clk);
#1;data_in = testData6[10491];
@(posedge clk);
#1;data_in = testData6[10492];
@(posedge clk);
#1;data_in = testData6[10493];
@(posedge clk);
#1;data_in = testData6[10494];
@(posedge clk);
#1;data_in = testData6[10495];
@(posedge clk);
#1;data_in = testData6[10496];
@(posedge clk);
#1;data_in = testData6[10497];
@(posedge clk);
#1;data_in = testData6[10498];
@(posedge clk);
#1;data_in = testData6[10499];
@(posedge clk);
#1;data_in = testData6[10500];
@(posedge clk);
#1;data_in = testData6[10501];
@(posedge clk);
#1;data_in = testData6[10502];
@(posedge clk);
#1;data_in = testData6[10503];
@(posedge clk);
#1;data_in = testData6[10504];
@(posedge clk);
#1;data_in = testData6[10505];
@(posedge clk);
#1;data_in = testData6[10506];
@(posedge clk);
#1;data_in = testData6[10507];
@(posedge clk);
#1;data_in = testData6[10508];
@(posedge clk);
#1;data_in = testData6[10509];
@(posedge clk);
#1;data_in = testData6[10510];
@(posedge clk);
#1;data_in = testData6[10511];
@(posedge clk);
#1;data_in = testData6[10512];
@(posedge clk);
#1;data_in = testData6[10513];
@(posedge clk);
#1;data_in = testData6[10514];
@(posedge clk);
#1;data_in = testData6[10515];
@(posedge clk);
#1;data_in = testData6[10516];
@(posedge clk);
#1;data_in = testData6[10517];
@(posedge clk);
#1;data_in = testData6[10518];
@(posedge clk);
#1;data_in = testData6[10519];
@(posedge clk);
#1;data_in = testData6[10520];
@(posedge clk);
#1;data_in = testData6[10521];
@(posedge clk);
#1;data_in = testData6[10522];
@(posedge clk);
#1;data_in = testData6[10523];
@(posedge clk);
#1;data_in = testData6[10524];
@(posedge clk);
#1;data_in = testData6[10525];
@(posedge clk);
#1;data_in = testData6[10526];
@(posedge clk);
#1;data_in = testData6[10527];
@(posedge clk);
#1;data_in = testData6[10528];
@(posedge clk);
#1;data_in = testData6[10529];
@(posedge clk);
#1;data_in = testData6[10530];
@(posedge clk);
#1;data_in = testData6[10531];
@(posedge clk);
#1;data_in = testData6[10532];
@(posedge clk);
#1;data_in = testData6[10533];
@(posedge clk);
#1;data_in = testData6[10534];
@(posedge clk);
#1;data_in = testData6[10535];
@(posedge clk);
#1;data_in = testData6[10536];
@(posedge clk);
#1;data_in = testData6[10537];
@(posedge clk);
#1;data_in = testData6[10538];
@(posedge clk);
#1;data_in = testData6[10539];
@(posedge clk);
#1;data_in = testData6[10540];
@(posedge clk);
#1;data_in = testData6[10541];
@(posedge clk);
#1;data_in = testData6[10542];
@(posedge clk);
#1;data_in = testData6[10543];
@(posedge clk);
#1;data_in = testData6[10544];
@(posedge clk);
#1;data_in = testData6[10545];
@(posedge clk);
#1;data_in = testData6[10546];
@(posedge clk);
#1;data_in = testData6[10547];
@(posedge clk);
#1;data_in = testData6[10548];
@(posedge clk);
#1;data_in = testData6[10549];
@(posedge clk);
#1;data_in = testData6[10550];
@(posedge clk);
#1;data_in = testData6[10551];
@(posedge clk);
#1;data_in = testData6[10552];
@(posedge clk);
#1;data_in = testData6[10553];
@(posedge clk);
#1;data_in = testData6[10554];
@(posedge clk);
#1;data_in = testData6[10555];
@(posedge clk);
#1;data_in = testData6[10556];
@(posedge clk);
#1;data_in = testData6[10557];
@(posedge clk);
#1;data_in = testData6[10558];
@(posedge clk);
#1;data_in = testData6[10559];
@(posedge clk);
#1;data_in = testData6[10560];
@(posedge clk);
#1;data_in = testData6[10561];
@(posedge clk);
#1;data_in = testData6[10562];
@(posedge clk);
#1;data_in = testData6[10563];
@(posedge clk);
#1;data_in = testData6[10564];
@(posedge clk);
#1;data_in = testData6[10565];
@(posedge clk);
#1;data_in = testData6[10566];
@(posedge clk);
#1;data_in = testData6[10567];
@(posedge clk);
#1;data_in = testData6[10568];
@(posedge clk);
#1;data_in = testData6[10569];
@(posedge clk);
#1;data_in = testData6[10570];
@(posedge clk);
#1;data_in = testData6[10571];
@(posedge clk);
#1;data_in = testData6[10572];
@(posedge clk);
#1;data_in = testData6[10573];
@(posedge clk);
#1;data_in = testData6[10574];
@(posedge clk);
#1;data_in = testData6[10575];
@(posedge clk);
#1;data_in = testData6[10576];
@(posedge clk);
#1;data_in = testData6[10577];
@(posedge clk);
#1;data_in = testData6[10578];
@(posedge clk);
#1;data_in = testData6[10579];
@(posedge clk);
#1;data_in = testData6[10580];
@(posedge clk);
#1;data_in = testData6[10581];
@(posedge clk);
#1;data_in = testData6[10582];
@(posedge clk);
#1;data_in = testData6[10583];
@(posedge clk);
#1;data_in = testData6[10584];
@(posedge clk);
#1;data_in = testData6[10585];
@(posedge clk);
#1;data_in = testData6[10586];
@(posedge clk);
#1;data_in = testData6[10587];
@(posedge clk);
#1;data_in = testData6[10588];
@(posedge clk);
#1;data_in = testData6[10589];
@(posedge clk);
#1;data_in = testData6[10590];
@(posedge clk);
#1;data_in = testData6[10591];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[10592]; 
@(posedge clk);
#1;data_in = testData6[10593];
@(posedge clk);
#1;data_in = testData6[10594];
@(posedge clk);
#1;data_in = testData6[10595];
@(posedge clk);
#1;data_in = testData6[10596];
@(posedge clk);
#1;data_in = testData6[10597];
@(posedge clk);
#1;data_in = testData6[10598];
@(posedge clk);
#1;data_in = testData6[10599];
@(posedge clk);
#1;data_in = testData6[10600];
@(posedge clk);
#1;data_in = testData6[10601];
@(posedge clk);
#1;data_in = testData6[10602];
@(posedge clk);
#1;data_in = testData6[10603];
@(posedge clk);
#1;data_in = testData6[10604];
@(posedge clk);
#1;data_in = testData6[10605];
@(posedge clk);
#1;data_in = testData6[10606];
@(posedge clk);
#1;data_in = testData6[10607];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[10608];
@(posedge clk);
#1;data_in = testData6[10609];
@(posedge clk);
#1;data_in = testData6[10610];
@(posedge clk);
#1;data_in = testData6[10611];
@(posedge clk);
#1;data_in = testData6[10612];
@(posedge clk);
#1;data_in = testData6[10613];
@(posedge clk);
#1;data_in = testData6[10614];
@(posedge clk);
#1;data_in = testData6[10615];
@(posedge clk);
#1;data_in = testData6[10616];
@(posedge clk);
#1;data_in = testData6[10617];
@(posedge clk);
#1;data_in = testData6[10618];
@(posedge clk);
#1;data_in = testData6[10619];
@(posedge clk);
#1;data_in = testData6[10620];
@(posedge clk);
#1;data_in = testData6[10621];
@(posedge clk);
#1;data_in = testData6[10622];
@(posedge clk);
#1;data_in = testData6[10623];
@(posedge clk);
#1;data_in = testData6[10624];
@(posedge clk);
#1;data_in = testData6[10625];
@(posedge clk);
#1;data_in = testData6[10626];
@(posedge clk);
#1;data_in = testData6[10627];
@(posedge clk);
#1;data_in = testData6[10628];
@(posedge clk);
#1;data_in = testData6[10629];
@(posedge clk);
#1;data_in = testData6[10630];
@(posedge clk);
#1;data_in = testData6[10631];
@(posedge clk);
#1;data_in = testData6[10632];
@(posedge clk);
#1;data_in = testData6[10633];
@(posedge clk);
#1;data_in = testData6[10634];
@(posedge clk);
#1;data_in = testData6[10635];
@(posedge clk);
#1;data_in = testData6[10636];
@(posedge clk);
#1;data_in = testData6[10637];
@(posedge clk);
#1;data_in = testData6[10638];
@(posedge clk);
#1;data_in = testData6[10639];
@(posedge clk);
#1;data_in = testData6[10640];
@(posedge clk);
#1;data_in = testData6[10641];
@(posedge clk);
#1;data_in = testData6[10642];
@(posedge clk);
#1;data_in = testData6[10643];
@(posedge clk);
#1;data_in = testData6[10644];
@(posedge clk);
#1;data_in = testData6[10645];
@(posedge clk);
#1;data_in = testData6[10646];
@(posedge clk);
#1;data_in = testData6[10647];
@(posedge clk);
#1;data_in = testData6[10648];
@(posedge clk);
#1;data_in = testData6[10649];
@(posedge clk);
#1;data_in = testData6[10650];
@(posedge clk);
#1;data_in = testData6[10651];
@(posedge clk);
#1;data_in = testData6[10652];
@(posedge clk);
#1;data_in = testData6[10653];
@(posedge clk);
#1;data_in = testData6[10654];
@(posedge clk);
#1;data_in = testData6[10655];
@(posedge clk);
#1;data_in = testData6[10656];
@(posedge clk);
#1;data_in = testData6[10657];
@(posedge clk);
#1;data_in = testData6[10658];
@(posedge clk);
#1;data_in = testData6[10659];
@(posedge clk);
#1;data_in = testData6[10660];
@(posedge clk);
#1;data_in = testData6[10661];
@(posedge clk);
#1;data_in = testData6[10662];
@(posedge clk);
#1;data_in = testData6[10663];
@(posedge clk);
#1;data_in = testData6[10664];
@(posedge clk);
#1;data_in = testData6[10665];
@(posedge clk);
#1;data_in = testData6[10666];
@(posedge clk);
#1;data_in = testData6[10667];
@(posedge clk);
#1;data_in = testData6[10668];
@(posedge clk);
#1;data_in = testData6[10669];
@(posedge clk);
#1;data_in = testData6[10670];
@(posedge clk);
#1;data_in = testData6[10671];
@(posedge clk);
#1;data_in = testData6[10672];
@(posedge clk);
#1;data_in = testData6[10673];
@(posedge clk);
#1;data_in = testData6[10674];
@(posedge clk);
#1;data_in = testData6[10675];
@(posedge clk);
#1;data_in = testData6[10676];
@(posedge clk);
#1;data_in = testData6[10677];
@(posedge clk);
#1;data_in = testData6[10678];
@(posedge clk);
#1;data_in = testData6[10679];
@(posedge clk);
#1;data_in = testData6[10680];
@(posedge clk);
#1;data_in = testData6[10681];
@(posedge clk);
#1;data_in = testData6[10682];
@(posedge clk);
#1;data_in = testData6[10683];
@(posedge clk);
#1;data_in = testData6[10684];
@(posedge clk);
#1;data_in = testData6[10685];
@(posedge clk);
#1;data_in = testData6[10686];
@(posedge clk);
#1;data_in = testData6[10687];
@(posedge clk);
#1;data_in = testData6[10688];
@(posedge clk);
#1;data_in = testData6[10689];
@(posedge clk);
#1;data_in = testData6[10690];
@(posedge clk);
#1;data_in = testData6[10691];
@(posedge clk);
#1;data_in = testData6[10692];
@(posedge clk);
#1;data_in = testData6[10693];
@(posedge clk);
#1;data_in = testData6[10694];
@(posedge clk);
#1;data_in = testData6[10695];
@(posedge clk);
#1;data_in = testData6[10696];
@(posedge clk);
#1;data_in = testData6[10697];
@(posedge clk);
#1;data_in = testData6[10698];
@(posedge clk);
#1;data_in = testData6[10699];
@(posedge clk);
#1;data_in = testData6[10700];
@(posedge clk);
#1;data_in = testData6[10701];
@(posedge clk);
#1;data_in = testData6[10702];
@(posedge clk);
#1;data_in = testData6[10703];
@(posedge clk);
#1;data_in = testData6[10704];
@(posedge clk);
#1;data_in = testData6[10705];
@(posedge clk);
#1;data_in = testData6[10706];
@(posedge clk);
#1;data_in = testData6[10707];
@(posedge clk);
#1;data_in = testData6[10708];
@(posedge clk);
#1;data_in = testData6[10709];
@(posedge clk);
#1;data_in = testData6[10710];
@(posedge clk);
#1;data_in = testData6[10711];
@(posedge clk);
#1;data_in = testData6[10712];
@(posedge clk);
#1;data_in = testData6[10713];
@(posedge clk);
#1;data_in = testData6[10714];
@(posedge clk);
#1;data_in = testData6[10715];
@(posedge clk);
#1;data_in = testData6[10716];
@(posedge clk);
#1;data_in = testData6[10717];
@(posedge clk);
#1;data_in = testData6[10718];
@(posedge clk);
#1;data_in = testData6[10719];
@(posedge clk);
#1;data_in = testData6[10720];
@(posedge clk);
#1;data_in = testData6[10721];
@(posedge clk);
#1;data_in = testData6[10722];
@(posedge clk);
#1;data_in = testData6[10723];
@(posedge clk);
#1;data_in = testData6[10724];
@(posedge clk);
#1;data_in = testData6[10725];
@(posedge clk);
#1;data_in = testData6[10726];
@(posedge clk);
#1;data_in = testData6[10727];
@(posedge clk);
#1;data_in = testData6[10728];
@(posedge clk);
#1;data_in = testData6[10729];
@(posedge clk);
#1;data_in = testData6[10730];
@(posedge clk);
#1;data_in = testData6[10731];
@(posedge clk);
#1;data_in = testData6[10732];
@(posedge clk);
#1;data_in = testData6[10733];
@(posedge clk);
#1;data_in = testData6[10734];
@(posedge clk);
#1;data_in = testData6[10735];
@(posedge clk);
#1;data_in = testData6[10736];
@(posedge clk);
#1;data_in = testData6[10737];
@(posedge clk);
#1;data_in = testData6[10738];
@(posedge clk);
#1;data_in = testData6[10739];
@(posedge clk);
#1;data_in = testData6[10740];
@(posedge clk);
#1;data_in = testData6[10741];
@(posedge clk);
#1;data_in = testData6[10742];
@(posedge clk);
#1;data_in = testData6[10743];
@(posedge clk);
#1;data_in = testData6[10744];
@(posedge clk);
#1;data_in = testData6[10745];
@(posedge clk);
#1;data_in = testData6[10746];
@(posedge clk);
#1;data_in = testData6[10747];
@(posedge clk);
#1;data_in = testData6[10748];
@(posedge clk);
#1;data_in = testData6[10749];
@(posedge clk);
#1;data_in = testData6[10750];
@(posedge clk);
#1;data_in = testData6[10751];
@(posedge clk);
#1;data_in = testData6[10752];
@(posedge clk);
#1;data_in = testData6[10753];
@(posedge clk);
#1;data_in = testData6[10754];
@(posedge clk);
#1;data_in = testData6[10755];
@(posedge clk);
#1;data_in = testData6[10756];
@(posedge clk);
#1;data_in = testData6[10757];
@(posedge clk);
#1;data_in = testData6[10758];
@(posedge clk);
#1;data_in = testData6[10759];
@(posedge clk);
#1;data_in = testData6[10760];
@(posedge clk);
#1;data_in = testData6[10761];
@(posedge clk);
#1;data_in = testData6[10762];
@(posedge clk);
#1;data_in = testData6[10763];
@(posedge clk);
#1;data_in = testData6[10764];
@(posedge clk);
#1;data_in = testData6[10765];
@(posedge clk);
#1;data_in = testData6[10766];
@(posedge clk);
#1;data_in = testData6[10767];
@(posedge clk);
#1;data_in = testData6[10768];
@(posedge clk);
#1;data_in = testData6[10769];
@(posedge clk);
#1;data_in = testData6[10770];
@(posedge clk);
#1;data_in = testData6[10771];
@(posedge clk);
#1;data_in = testData6[10772];
@(posedge clk);
#1;data_in = testData6[10773];
@(posedge clk);
#1;data_in = testData6[10774];
@(posedge clk);
#1;data_in = testData6[10775];
@(posedge clk);
#1;data_in = testData6[10776];
@(posedge clk);
#1;data_in = testData6[10777];
@(posedge clk);
#1;data_in = testData6[10778];
@(posedge clk);
#1;data_in = testData6[10779];
@(posedge clk);
#1;data_in = testData6[10780];
@(posedge clk);
#1;data_in = testData6[10781];
@(posedge clk);
#1;data_in = testData6[10782];
@(posedge clk);
#1;data_in = testData6[10783];
@(posedge clk);
#1;data_in = testData6[10784];
@(posedge clk);
#1;data_in = testData6[10785];
@(posedge clk);
#1;data_in = testData6[10786];
@(posedge clk);
#1;data_in = testData6[10787];
@(posedge clk);
#1;data_in = testData6[10788];
@(posedge clk);
#1;data_in = testData6[10789];
@(posedge clk);
#1;data_in = testData6[10790];
@(posedge clk);
#1;data_in = testData6[10791];
@(posedge clk);
#1;data_in = testData6[10792];
@(posedge clk);
#1;data_in = testData6[10793];
@(posedge clk);
#1;data_in = testData6[10794];
@(posedge clk);
#1;data_in = testData6[10795];
@(posedge clk);
#1;data_in = testData6[10796];
@(posedge clk);
#1;data_in = testData6[10797];
@(posedge clk);
#1;data_in = testData6[10798];
@(posedge clk);
#1;data_in = testData6[10799];
@(posedge clk);
#1;data_in = testData6[10800];
@(posedge clk);
#1;data_in = testData6[10801];
@(posedge clk);
#1;data_in = testData6[10802];
@(posedge clk);
#1;data_in = testData6[10803];
@(posedge clk);
#1;data_in = testData6[10804];
@(posedge clk);
#1;data_in = testData6[10805];
@(posedge clk);
#1;data_in = testData6[10806];
@(posedge clk);
#1;data_in = testData6[10807];
@(posedge clk);
#1;data_in = testData6[10808];
@(posedge clk);
#1;data_in = testData6[10809];
@(posedge clk);
#1;data_in = testData6[10810];
@(posedge clk);
#1;data_in = testData6[10811];
@(posedge clk);
#1;data_in = testData6[10812];
@(posedge clk);
#1;data_in = testData6[10813];
@(posedge clk);
#1;data_in = testData6[10814];
@(posedge clk);
#1;data_in = testData6[10815];
@(posedge clk);
#1;data_in = testData6[10816];
@(posedge clk);
#1;data_in = testData6[10817];
@(posedge clk);
#1;data_in = testData6[10818];
@(posedge clk);
#1;data_in = testData6[10819];
@(posedge clk);
#1;data_in = testData6[10820];
@(posedge clk);
#1;data_in = testData6[10821];
@(posedge clk);
#1;data_in = testData6[10822];
@(posedge clk);
#1;data_in = testData6[10823];
@(posedge clk);
#1;data_in = testData6[10824];
@(posedge clk);
#1;data_in = testData6[10825];
@(posedge clk);
#1;data_in = testData6[10826];
@(posedge clk);
#1;data_in = testData6[10827];
@(posedge clk);
#1;data_in = testData6[10828];
@(posedge clk);
#1;data_in = testData6[10829];
@(posedge clk);
#1;data_in = testData6[10830];
@(posedge clk);
#1;data_in = testData6[10831];
@(posedge clk);
#1;data_in = testData6[10832];
@(posedge clk);
#1;data_in = testData6[10833];
@(posedge clk);
#1;data_in = testData6[10834];
@(posedge clk);
#1;data_in = testData6[10835];
@(posedge clk);
#1;data_in = testData6[10836];
@(posedge clk);
#1;data_in = testData6[10837];
@(posedge clk);
#1;data_in = testData6[10838];
@(posedge clk);
#1;data_in = testData6[10839];
@(posedge clk);
#1;data_in = testData6[10840];
@(posedge clk);
#1;data_in = testData6[10841];
@(posedge clk);
#1;data_in = testData6[10842];
@(posedge clk);
#1;data_in = testData6[10843];
@(posedge clk);
#1;data_in = testData6[10844];
@(posedge clk);
#1;data_in = testData6[10845];
@(posedge clk);
#1;data_in = testData6[10846];
@(posedge clk);
#1;data_in = testData6[10847];
@(posedge clk);
#1;data_in = testData6[10848];
@(posedge clk);
#1;data_in = testData6[10849];
@(posedge clk);
#1;data_in = testData6[10850];
@(posedge clk);
#1;data_in = testData6[10851];
@(posedge clk);
#1;data_in = testData6[10852];
@(posedge clk);
#1;data_in = testData6[10853];
@(posedge clk);
#1;data_in = testData6[10854];
@(posedge clk);
#1;data_in = testData6[10855];
@(posedge clk);
#1;data_in = testData6[10856];
@(posedge clk);
#1;data_in = testData6[10857];
@(posedge clk);
#1;data_in = testData6[10858];
@(posedge clk);
#1;data_in = testData6[10859];
@(posedge clk);
#1;data_in = testData6[10860];
@(posedge clk);
#1;data_in = testData6[10861];
@(posedge clk);
#1;data_in = testData6[10862];
@(posedge clk);
#1;data_in = testData6[10863];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[10864]; 
@(posedge clk);
#1;data_in = testData6[10865];
@(posedge clk);
#1;data_in = testData6[10866];
@(posedge clk);
#1;data_in = testData6[10867];
@(posedge clk);
#1;data_in = testData6[10868];
@(posedge clk);
#1;data_in = testData6[10869];
@(posedge clk);
#1;data_in = testData6[10870];
@(posedge clk);
#1;data_in = testData6[10871];
@(posedge clk);
#1;data_in = testData6[10872];
@(posedge clk);
#1;data_in = testData6[10873];
@(posedge clk);
#1;data_in = testData6[10874];
@(posedge clk);
#1;data_in = testData6[10875];
@(posedge clk);
#1;data_in = testData6[10876];
@(posedge clk);
#1;data_in = testData6[10877];
@(posedge clk);
#1;data_in = testData6[10878];
@(posedge clk);
#1;data_in = testData6[10879];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[10880];
@(posedge clk);
#1;data_in = testData6[10881];
@(posedge clk);
#1;data_in = testData6[10882];
@(posedge clk);
#1;data_in = testData6[10883];
@(posedge clk);
#1;data_in = testData6[10884];
@(posedge clk);
#1;data_in = testData6[10885];
@(posedge clk);
#1;data_in = testData6[10886];
@(posedge clk);
#1;data_in = testData6[10887];
@(posedge clk);
#1;data_in = testData6[10888];
@(posedge clk);
#1;data_in = testData6[10889];
@(posedge clk);
#1;data_in = testData6[10890];
@(posedge clk);
#1;data_in = testData6[10891];
@(posedge clk);
#1;data_in = testData6[10892];
@(posedge clk);
#1;data_in = testData6[10893];
@(posedge clk);
#1;data_in = testData6[10894];
@(posedge clk);
#1;data_in = testData6[10895];
@(posedge clk);
#1;data_in = testData6[10896];
@(posedge clk);
#1;data_in = testData6[10897];
@(posedge clk);
#1;data_in = testData6[10898];
@(posedge clk);
#1;data_in = testData6[10899];
@(posedge clk);
#1;data_in = testData6[10900];
@(posedge clk);
#1;data_in = testData6[10901];
@(posedge clk);
#1;data_in = testData6[10902];
@(posedge clk);
#1;data_in = testData6[10903];
@(posedge clk);
#1;data_in = testData6[10904];
@(posedge clk);
#1;data_in = testData6[10905];
@(posedge clk);
#1;data_in = testData6[10906];
@(posedge clk);
#1;data_in = testData6[10907];
@(posedge clk);
#1;data_in = testData6[10908];
@(posedge clk);
#1;data_in = testData6[10909];
@(posedge clk);
#1;data_in = testData6[10910];
@(posedge clk);
#1;data_in = testData6[10911];
@(posedge clk);
#1;data_in = testData6[10912];
@(posedge clk);
#1;data_in = testData6[10913];
@(posedge clk);
#1;data_in = testData6[10914];
@(posedge clk);
#1;data_in = testData6[10915];
@(posedge clk);
#1;data_in = testData6[10916];
@(posedge clk);
#1;data_in = testData6[10917];
@(posedge clk);
#1;data_in = testData6[10918];
@(posedge clk);
#1;data_in = testData6[10919];
@(posedge clk);
#1;data_in = testData6[10920];
@(posedge clk);
#1;data_in = testData6[10921];
@(posedge clk);
#1;data_in = testData6[10922];
@(posedge clk);
#1;data_in = testData6[10923];
@(posedge clk);
#1;data_in = testData6[10924];
@(posedge clk);
#1;data_in = testData6[10925];
@(posedge clk);
#1;data_in = testData6[10926];
@(posedge clk);
#1;data_in = testData6[10927];
@(posedge clk);
#1;data_in = testData6[10928];
@(posedge clk);
#1;data_in = testData6[10929];
@(posedge clk);
#1;data_in = testData6[10930];
@(posedge clk);
#1;data_in = testData6[10931];
@(posedge clk);
#1;data_in = testData6[10932];
@(posedge clk);
#1;data_in = testData6[10933];
@(posedge clk);
#1;data_in = testData6[10934];
@(posedge clk);
#1;data_in = testData6[10935];
@(posedge clk);
#1;data_in = testData6[10936];
@(posedge clk);
#1;data_in = testData6[10937];
@(posedge clk);
#1;data_in = testData6[10938];
@(posedge clk);
#1;data_in = testData6[10939];
@(posedge clk);
#1;data_in = testData6[10940];
@(posedge clk);
#1;data_in = testData6[10941];
@(posedge clk);
#1;data_in = testData6[10942];
@(posedge clk);
#1;data_in = testData6[10943];
@(posedge clk);
#1;data_in = testData6[10944];
@(posedge clk);
#1;data_in = testData6[10945];
@(posedge clk);
#1;data_in = testData6[10946];
@(posedge clk);
#1;data_in = testData6[10947];
@(posedge clk);
#1;data_in = testData6[10948];
@(posedge clk);
#1;data_in = testData6[10949];
@(posedge clk);
#1;data_in = testData6[10950];
@(posedge clk);
#1;data_in = testData6[10951];
@(posedge clk);
#1;data_in = testData6[10952];
@(posedge clk);
#1;data_in = testData6[10953];
@(posedge clk);
#1;data_in = testData6[10954];
@(posedge clk);
#1;data_in = testData6[10955];
@(posedge clk);
#1;data_in = testData6[10956];
@(posedge clk);
#1;data_in = testData6[10957];
@(posedge clk);
#1;data_in = testData6[10958];
@(posedge clk);
#1;data_in = testData6[10959];
@(posedge clk);
#1;data_in = testData6[10960];
@(posedge clk);
#1;data_in = testData6[10961];
@(posedge clk);
#1;data_in = testData6[10962];
@(posedge clk);
#1;data_in = testData6[10963];
@(posedge clk);
#1;data_in = testData6[10964];
@(posedge clk);
#1;data_in = testData6[10965];
@(posedge clk);
#1;data_in = testData6[10966];
@(posedge clk);
#1;data_in = testData6[10967];
@(posedge clk);
#1;data_in = testData6[10968];
@(posedge clk);
#1;data_in = testData6[10969];
@(posedge clk);
#1;data_in = testData6[10970];
@(posedge clk);
#1;data_in = testData6[10971];
@(posedge clk);
#1;data_in = testData6[10972];
@(posedge clk);
#1;data_in = testData6[10973];
@(posedge clk);
#1;data_in = testData6[10974];
@(posedge clk);
#1;data_in = testData6[10975];
@(posedge clk);
#1;data_in = testData6[10976];
@(posedge clk);
#1;data_in = testData6[10977];
@(posedge clk);
#1;data_in = testData6[10978];
@(posedge clk);
#1;data_in = testData6[10979];
@(posedge clk);
#1;data_in = testData6[10980];
@(posedge clk);
#1;data_in = testData6[10981];
@(posedge clk);
#1;data_in = testData6[10982];
@(posedge clk);
#1;data_in = testData6[10983];
@(posedge clk);
#1;data_in = testData6[10984];
@(posedge clk);
#1;data_in = testData6[10985];
@(posedge clk);
#1;data_in = testData6[10986];
@(posedge clk);
#1;data_in = testData6[10987];
@(posedge clk);
#1;data_in = testData6[10988];
@(posedge clk);
#1;data_in = testData6[10989];
@(posedge clk);
#1;data_in = testData6[10990];
@(posedge clk);
#1;data_in = testData6[10991];
@(posedge clk);
#1;data_in = testData6[10992];
@(posedge clk);
#1;data_in = testData6[10993];
@(posedge clk);
#1;data_in = testData6[10994];
@(posedge clk);
#1;data_in = testData6[10995];
@(posedge clk);
#1;data_in = testData6[10996];
@(posedge clk);
#1;data_in = testData6[10997];
@(posedge clk);
#1;data_in = testData6[10998];
@(posedge clk);
#1;data_in = testData6[10999];
@(posedge clk);
#1;data_in = testData6[11000];
@(posedge clk);
#1;data_in = testData6[11001];
@(posedge clk);
#1;data_in = testData6[11002];
@(posedge clk);
#1;data_in = testData6[11003];
@(posedge clk);
#1;data_in = testData6[11004];
@(posedge clk);
#1;data_in = testData6[11005];
@(posedge clk);
#1;data_in = testData6[11006];
@(posedge clk);
#1;data_in = testData6[11007];
@(posedge clk);
#1;data_in = testData6[11008];
@(posedge clk);
#1;data_in = testData6[11009];
@(posedge clk);
#1;data_in = testData6[11010];
@(posedge clk);
#1;data_in = testData6[11011];
@(posedge clk);
#1;data_in = testData6[11012];
@(posedge clk);
#1;data_in = testData6[11013];
@(posedge clk);
#1;data_in = testData6[11014];
@(posedge clk);
#1;data_in = testData6[11015];
@(posedge clk);
#1;data_in = testData6[11016];
@(posedge clk);
#1;data_in = testData6[11017];
@(posedge clk);
#1;data_in = testData6[11018];
@(posedge clk);
#1;data_in = testData6[11019];
@(posedge clk);
#1;data_in = testData6[11020];
@(posedge clk);
#1;data_in = testData6[11021];
@(posedge clk);
#1;data_in = testData6[11022];
@(posedge clk);
#1;data_in = testData6[11023];
@(posedge clk);
#1;data_in = testData6[11024];
@(posedge clk);
#1;data_in = testData6[11025];
@(posedge clk);
#1;data_in = testData6[11026];
@(posedge clk);
#1;data_in = testData6[11027];
@(posedge clk);
#1;data_in = testData6[11028];
@(posedge clk);
#1;data_in = testData6[11029];
@(posedge clk);
#1;data_in = testData6[11030];
@(posedge clk);
#1;data_in = testData6[11031];
@(posedge clk);
#1;data_in = testData6[11032];
@(posedge clk);
#1;data_in = testData6[11033];
@(posedge clk);
#1;data_in = testData6[11034];
@(posedge clk);
#1;data_in = testData6[11035];
@(posedge clk);
#1;data_in = testData6[11036];
@(posedge clk);
#1;data_in = testData6[11037];
@(posedge clk);
#1;data_in = testData6[11038];
@(posedge clk);
#1;data_in = testData6[11039];
@(posedge clk);
#1;data_in = testData6[11040];
@(posedge clk);
#1;data_in = testData6[11041];
@(posedge clk);
#1;data_in = testData6[11042];
@(posedge clk);
#1;data_in = testData6[11043];
@(posedge clk);
#1;data_in = testData6[11044];
@(posedge clk);
#1;data_in = testData6[11045];
@(posedge clk);
#1;data_in = testData6[11046];
@(posedge clk);
#1;data_in = testData6[11047];
@(posedge clk);
#1;data_in = testData6[11048];
@(posedge clk);
#1;data_in = testData6[11049];
@(posedge clk);
#1;data_in = testData6[11050];
@(posedge clk);
#1;data_in = testData6[11051];
@(posedge clk);
#1;data_in = testData6[11052];
@(posedge clk);
#1;data_in = testData6[11053];
@(posedge clk);
#1;data_in = testData6[11054];
@(posedge clk);
#1;data_in = testData6[11055];
@(posedge clk);
#1;data_in = testData6[11056];
@(posedge clk);
#1;data_in = testData6[11057];
@(posedge clk);
#1;data_in = testData6[11058];
@(posedge clk);
#1;data_in = testData6[11059];
@(posedge clk);
#1;data_in = testData6[11060];
@(posedge clk);
#1;data_in = testData6[11061];
@(posedge clk);
#1;data_in = testData6[11062];
@(posedge clk);
#1;data_in = testData6[11063];
@(posedge clk);
#1;data_in = testData6[11064];
@(posedge clk);
#1;data_in = testData6[11065];
@(posedge clk);
#1;data_in = testData6[11066];
@(posedge clk);
#1;data_in = testData6[11067];
@(posedge clk);
#1;data_in = testData6[11068];
@(posedge clk);
#1;data_in = testData6[11069];
@(posedge clk);
#1;data_in = testData6[11070];
@(posedge clk);
#1;data_in = testData6[11071];
@(posedge clk);
#1;data_in = testData6[11072];
@(posedge clk);
#1;data_in = testData6[11073];
@(posedge clk);
#1;data_in = testData6[11074];
@(posedge clk);
#1;data_in = testData6[11075];
@(posedge clk);
#1;data_in = testData6[11076];
@(posedge clk);
#1;data_in = testData6[11077];
@(posedge clk);
#1;data_in = testData6[11078];
@(posedge clk);
#1;data_in = testData6[11079];
@(posedge clk);
#1;data_in = testData6[11080];
@(posedge clk);
#1;data_in = testData6[11081];
@(posedge clk);
#1;data_in = testData6[11082];
@(posedge clk);
#1;data_in = testData6[11083];
@(posedge clk);
#1;data_in = testData6[11084];
@(posedge clk);
#1;data_in = testData6[11085];
@(posedge clk);
#1;data_in = testData6[11086];
@(posedge clk);
#1;data_in = testData6[11087];
@(posedge clk);
#1;data_in = testData6[11088];
@(posedge clk);
#1;data_in = testData6[11089];
@(posedge clk);
#1;data_in = testData6[11090];
@(posedge clk);
#1;data_in = testData6[11091];
@(posedge clk);
#1;data_in = testData6[11092];
@(posedge clk);
#1;data_in = testData6[11093];
@(posedge clk);
#1;data_in = testData6[11094];
@(posedge clk);
#1;data_in = testData6[11095];
@(posedge clk);
#1;data_in = testData6[11096];
@(posedge clk);
#1;data_in = testData6[11097];
@(posedge clk);
#1;data_in = testData6[11098];
@(posedge clk);
#1;data_in = testData6[11099];
@(posedge clk);
#1;data_in = testData6[11100];
@(posedge clk);
#1;data_in = testData6[11101];
@(posedge clk);
#1;data_in = testData6[11102];
@(posedge clk);
#1;data_in = testData6[11103];
@(posedge clk);
#1;data_in = testData6[11104];
@(posedge clk);
#1;data_in = testData6[11105];
@(posedge clk);
#1;data_in = testData6[11106];
@(posedge clk);
#1;data_in = testData6[11107];
@(posedge clk);
#1;data_in = testData6[11108];
@(posedge clk);
#1;data_in = testData6[11109];
@(posedge clk);
#1;data_in = testData6[11110];
@(posedge clk);
#1;data_in = testData6[11111];
@(posedge clk);
#1;data_in = testData6[11112];
@(posedge clk);
#1;data_in = testData6[11113];
@(posedge clk);
#1;data_in = testData6[11114];
@(posedge clk);
#1;data_in = testData6[11115];
@(posedge clk);
#1;data_in = testData6[11116];
@(posedge clk);
#1;data_in = testData6[11117];
@(posedge clk);
#1;data_in = testData6[11118];
@(posedge clk);
#1;data_in = testData6[11119];
@(posedge clk);
#1;data_in = testData6[11120];
@(posedge clk);
#1;data_in = testData6[11121];
@(posedge clk);
#1;data_in = testData6[11122];
@(posedge clk);
#1;data_in = testData6[11123];
@(posedge clk);
#1;data_in = testData6[11124];
@(posedge clk);
#1;data_in = testData6[11125];
@(posedge clk);
#1;data_in = testData6[11126];
@(posedge clk);
#1;data_in = testData6[11127];
@(posedge clk);
#1;data_in = testData6[11128];
@(posedge clk);
#1;data_in = testData6[11129];
@(posedge clk);
#1;data_in = testData6[11130];
@(posedge clk);
#1;data_in = testData6[11131];
@(posedge clk);
#1;data_in = testData6[11132];
@(posedge clk);
#1;data_in = testData6[11133];
@(posedge clk);
#1;data_in = testData6[11134];
@(posedge clk);
#1;data_in = testData6[11135];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[11136]; 
@(posedge clk);
#1;data_in = testData6[11137];
@(posedge clk);
#1;data_in = testData6[11138];
@(posedge clk);
#1;data_in = testData6[11139];
@(posedge clk);
#1;data_in = testData6[11140];
@(posedge clk);
#1;data_in = testData6[11141];
@(posedge clk);
#1;data_in = testData6[11142];
@(posedge clk);
#1;data_in = testData6[11143];
@(posedge clk);
#1;data_in = testData6[11144];
@(posedge clk);
#1;data_in = testData6[11145];
@(posedge clk);
#1;data_in = testData6[11146];
@(posedge clk);
#1;data_in = testData6[11147];
@(posedge clk);
#1;data_in = testData6[11148];
@(posedge clk);
#1;data_in = testData6[11149];
@(posedge clk);
#1;data_in = testData6[11150];
@(posedge clk);
#1;data_in = testData6[11151];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[11152];
@(posedge clk);
#1;data_in = testData6[11153];
@(posedge clk);
#1;data_in = testData6[11154];
@(posedge clk);
#1;data_in = testData6[11155];
@(posedge clk);
#1;data_in = testData6[11156];
@(posedge clk);
#1;data_in = testData6[11157];
@(posedge clk);
#1;data_in = testData6[11158];
@(posedge clk);
#1;data_in = testData6[11159];
@(posedge clk);
#1;data_in = testData6[11160];
@(posedge clk);
#1;data_in = testData6[11161];
@(posedge clk);
#1;data_in = testData6[11162];
@(posedge clk);
#1;data_in = testData6[11163];
@(posedge clk);
#1;data_in = testData6[11164];
@(posedge clk);
#1;data_in = testData6[11165];
@(posedge clk);
#1;data_in = testData6[11166];
@(posedge clk);
#1;data_in = testData6[11167];
@(posedge clk);
#1;data_in = testData6[11168];
@(posedge clk);
#1;data_in = testData6[11169];
@(posedge clk);
#1;data_in = testData6[11170];
@(posedge clk);
#1;data_in = testData6[11171];
@(posedge clk);
#1;data_in = testData6[11172];
@(posedge clk);
#1;data_in = testData6[11173];
@(posedge clk);
#1;data_in = testData6[11174];
@(posedge clk);
#1;data_in = testData6[11175];
@(posedge clk);
#1;data_in = testData6[11176];
@(posedge clk);
#1;data_in = testData6[11177];
@(posedge clk);
#1;data_in = testData6[11178];
@(posedge clk);
#1;data_in = testData6[11179];
@(posedge clk);
#1;data_in = testData6[11180];
@(posedge clk);
#1;data_in = testData6[11181];
@(posedge clk);
#1;data_in = testData6[11182];
@(posedge clk);
#1;data_in = testData6[11183];
@(posedge clk);
#1;data_in = testData6[11184];
@(posedge clk);
#1;data_in = testData6[11185];
@(posedge clk);
#1;data_in = testData6[11186];
@(posedge clk);
#1;data_in = testData6[11187];
@(posedge clk);
#1;data_in = testData6[11188];
@(posedge clk);
#1;data_in = testData6[11189];
@(posedge clk);
#1;data_in = testData6[11190];
@(posedge clk);
#1;data_in = testData6[11191];
@(posedge clk);
#1;data_in = testData6[11192];
@(posedge clk);
#1;data_in = testData6[11193];
@(posedge clk);
#1;data_in = testData6[11194];
@(posedge clk);
#1;data_in = testData6[11195];
@(posedge clk);
#1;data_in = testData6[11196];
@(posedge clk);
#1;data_in = testData6[11197];
@(posedge clk);
#1;data_in = testData6[11198];
@(posedge clk);
#1;data_in = testData6[11199];
@(posedge clk);
#1;data_in = testData6[11200];
@(posedge clk);
#1;data_in = testData6[11201];
@(posedge clk);
#1;data_in = testData6[11202];
@(posedge clk);
#1;data_in = testData6[11203];
@(posedge clk);
#1;data_in = testData6[11204];
@(posedge clk);
#1;data_in = testData6[11205];
@(posedge clk);
#1;data_in = testData6[11206];
@(posedge clk);
#1;data_in = testData6[11207];
@(posedge clk);
#1;data_in = testData6[11208];
@(posedge clk);
#1;data_in = testData6[11209];
@(posedge clk);
#1;data_in = testData6[11210];
@(posedge clk);
#1;data_in = testData6[11211];
@(posedge clk);
#1;data_in = testData6[11212];
@(posedge clk);
#1;data_in = testData6[11213];
@(posedge clk);
#1;data_in = testData6[11214];
@(posedge clk);
#1;data_in = testData6[11215];
@(posedge clk);
#1;data_in = testData6[11216];
@(posedge clk);
#1;data_in = testData6[11217];
@(posedge clk);
#1;data_in = testData6[11218];
@(posedge clk);
#1;data_in = testData6[11219];
@(posedge clk);
#1;data_in = testData6[11220];
@(posedge clk);
#1;data_in = testData6[11221];
@(posedge clk);
#1;data_in = testData6[11222];
@(posedge clk);
#1;data_in = testData6[11223];
@(posedge clk);
#1;data_in = testData6[11224];
@(posedge clk);
#1;data_in = testData6[11225];
@(posedge clk);
#1;data_in = testData6[11226];
@(posedge clk);
#1;data_in = testData6[11227];
@(posedge clk);
#1;data_in = testData6[11228];
@(posedge clk);
#1;data_in = testData6[11229];
@(posedge clk);
#1;data_in = testData6[11230];
@(posedge clk);
#1;data_in = testData6[11231];
@(posedge clk);
#1;data_in = testData6[11232];
@(posedge clk);
#1;data_in = testData6[11233];
@(posedge clk);
#1;data_in = testData6[11234];
@(posedge clk);
#1;data_in = testData6[11235];
@(posedge clk);
#1;data_in = testData6[11236];
@(posedge clk);
#1;data_in = testData6[11237];
@(posedge clk);
#1;data_in = testData6[11238];
@(posedge clk);
#1;data_in = testData6[11239];
@(posedge clk);
#1;data_in = testData6[11240];
@(posedge clk);
#1;data_in = testData6[11241];
@(posedge clk);
#1;data_in = testData6[11242];
@(posedge clk);
#1;data_in = testData6[11243];
@(posedge clk);
#1;data_in = testData6[11244];
@(posedge clk);
#1;data_in = testData6[11245];
@(posedge clk);
#1;data_in = testData6[11246];
@(posedge clk);
#1;data_in = testData6[11247];
@(posedge clk);
#1;data_in = testData6[11248];
@(posedge clk);
#1;data_in = testData6[11249];
@(posedge clk);
#1;data_in = testData6[11250];
@(posedge clk);
#1;data_in = testData6[11251];
@(posedge clk);
#1;data_in = testData6[11252];
@(posedge clk);
#1;data_in = testData6[11253];
@(posedge clk);
#1;data_in = testData6[11254];
@(posedge clk);
#1;data_in = testData6[11255];
@(posedge clk);
#1;data_in = testData6[11256];
@(posedge clk);
#1;data_in = testData6[11257];
@(posedge clk);
#1;data_in = testData6[11258];
@(posedge clk);
#1;data_in = testData6[11259];
@(posedge clk);
#1;data_in = testData6[11260];
@(posedge clk);
#1;data_in = testData6[11261];
@(posedge clk);
#1;data_in = testData6[11262];
@(posedge clk);
#1;data_in = testData6[11263];
@(posedge clk);
#1;data_in = testData6[11264];
@(posedge clk);
#1;data_in = testData6[11265];
@(posedge clk);
#1;data_in = testData6[11266];
@(posedge clk);
#1;data_in = testData6[11267];
@(posedge clk);
#1;data_in = testData6[11268];
@(posedge clk);
#1;data_in = testData6[11269];
@(posedge clk);
#1;data_in = testData6[11270];
@(posedge clk);
#1;data_in = testData6[11271];
@(posedge clk);
#1;data_in = testData6[11272];
@(posedge clk);
#1;data_in = testData6[11273];
@(posedge clk);
#1;data_in = testData6[11274];
@(posedge clk);
#1;data_in = testData6[11275];
@(posedge clk);
#1;data_in = testData6[11276];
@(posedge clk);
#1;data_in = testData6[11277];
@(posedge clk);
#1;data_in = testData6[11278];
@(posedge clk);
#1;data_in = testData6[11279];
@(posedge clk);
#1;data_in = testData6[11280];
@(posedge clk);
#1;data_in = testData6[11281];
@(posedge clk);
#1;data_in = testData6[11282];
@(posedge clk);
#1;data_in = testData6[11283];
@(posedge clk);
#1;data_in = testData6[11284];
@(posedge clk);
#1;data_in = testData6[11285];
@(posedge clk);
#1;data_in = testData6[11286];
@(posedge clk);
#1;data_in = testData6[11287];
@(posedge clk);
#1;data_in = testData6[11288];
@(posedge clk);
#1;data_in = testData6[11289];
@(posedge clk);
#1;data_in = testData6[11290];
@(posedge clk);
#1;data_in = testData6[11291];
@(posedge clk);
#1;data_in = testData6[11292];
@(posedge clk);
#1;data_in = testData6[11293];
@(posedge clk);
#1;data_in = testData6[11294];
@(posedge clk);
#1;data_in = testData6[11295];
@(posedge clk);
#1;data_in = testData6[11296];
@(posedge clk);
#1;data_in = testData6[11297];
@(posedge clk);
#1;data_in = testData6[11298];
@(posedge clk);
#1;data_in = testData6[11299];
@(posedge clk);
#1;data_in = testData6[11300];
@(posedge clk);
#1;data_in = testData6[11301];
@(posedge clk);
#1;data_in = testData6[11302];
@(posedge clk);
#1;data_in = testData6[11303];
@(posedge clk);
#1;data_in = testData6[11304];
@(posedge clk);
#1;data_in = testData6[11305];
@(posedge clk);
#1;data_in = testData6[11306];
@(posedge clk);
#1;data_in = testData6[11307];
@(posedge clk);
#1;data_in = testData6[11308];
@(posedge clk);
#1;data_in = testData6[11309];
@(posedge clk);
#1;data_in = testData6[11310];
@(posedge clk);
#1;data_in = testData6[11311];
@(posedge clk);
#1;data_in = testData6[11312];
@(posedge clk);
#1;data_in = testData6[11313];
@(posedge clk);
#1;data_in = testData6[11314];
@(posedge clk);
#1;data_in = testData6[11315];
@(posedge clk);
#1;data_in = testData6[11316];
@(posedge clk);
#1;data_in = testData6[11317];
@(posedge clk);
#1;data_in = testData6[11318];
@(posedge clk);
#1;data_in = testData6[11319];
@(posedge clk);
#1;data_in = testData6[11320];
@(posedge clk);
#1;data_in = testData6[11321];
@(posedge clk);
#1;data_in = testData6[11322];
@(posedge clk);
#1;data_in = testData6[11323];
@(posedge clk);
#1;data_in = testData6[11324];
@(posedge clk);
#1;data_in = testData6[11325];
@(posedge clk);
#1;data_in = testData6[11326];
@(posedge clk);
#1;data_in = testData6[11327];
@(posedge clk);
#1;data_in = testData6[11328];
@(posedge clk);
#1;data_in = testData6[11329];
@(posedge clk);
#1;data_in = testData6[11330];
@(posedge clk);
#1;data_in = testData6[11331];
@(posedge clk);
#1;data_in = testData6[11332];
@(posedge clk);
#1;data_in = testData6[11333];
@(posedge clk);
#1;data_in = testData6[11334];
@(posedge clk);
#1;data_in = testData6[11335];
@(posedge clk);
#1;data_in = testData6[11336];
@(posedge clk);
#1;data_in = testData6[11337];
@(posedge clk);
#1;data_in = testData6[11338];
@(posedge clk);
#1;data_in = testData6[11339];
@(posedge clk);
#1;data_in = testData6[11340];
@(posedge clk);
#1;data_in = testData6[11341];
@(posedge clk);
#1;data_in = testData6[11342];
@(posedge clk);
#1;data_in = testData6[11343];
@(posedge clk);
#1;data_in = testData6[11344];
@(posedge clk);
#1;data_in = testData6[11345];
@(posedge clk);
#1;data_in = testData6[11346];
@(posedge clk);
#1;data_in = testData6[11347];
@(posedge clk);
#1;data_in = testData6[11348];
@(posedge clk);
#1;data_in = testData6[11349];
@(posedge clk);
#1;data_in = testData6[11350];
@(posedge clk);
#1;data_in = testData6[11351];
@(posedge clk);
#1;data_in = testData6[11352];
@(posedge clk);
#1;data_in = testData6[11353];
@(posedge clk);
#1;data_in = testData6[11354];
@(posedge clk);
#1;data_in = testData6[11355];
@(posedge clk);
#1;data_in = testData6[11356];
@(posedge clk);
#1;data_in = testData6[11357];
@(posedge clk);
#1;data_in = testData6[11358];
@(posedge clk);
#1;data_in = testData6[11359];
@(posedge clk);
#1;data_in = testData6[11360];
@(posedge clk);
#1;data_in = testData6[11361];
@(posedge clk);
#1;data_in = testData6[11362];
@(posedge clk);
#1;data_in = testData6[11363];
@(posedge clk);
#1;data_in = testData6[11364];
@(posedge clk);
#1;data_in = testData6[11365];
@(posedge clk);
#1;data_in = testData6[11366];
@(posedge clk);
#1;data_in = testData6[11367];
@(posedge clk);
#1;data_in = testData6[11368];
@(posedge clk);
#1;data_in = testData6[11369];
@(posedge clk);
#1;data_in = testData6[11370];
@(posedge clk);
#1;data_in = testData6[11371];
@(posedge clk);
#1;data_in = testData6[11372];
@(posedge clk);
#1;data_in = testData6[11373];
@(posedge clk);
#1;data_in = testData6[11374];
@(posedge clk);
#1;data_in = testData6[11375];
@(posedge clk);
#1;data_in = testData6[11376];
@(posedge clk);
#1;data_in = testData6[11377];
@(posedge clk);
#1;data_in = testData6[11378];
@(posedge clk);
#1;data_in = testData6[11379];
@(posedge clk);
#1;data_in = testData6[11380];
@(posedge clk);
#1;data_in = testData6[11381];
@(posedge clk);
#1;data_in = testData6[11382];
@(posedge clk);
#1;data_in = testData6[11383];
@(posedge clk);
#1;data_in = testData6[11384];
@(posedge clk);
#1;data_in = testData6[11385];
@(posedge clk);
#1;data_in = testData6[11386];
@(posedge clk);
#1;data_in = testData6[11387];
@(posedge clk);
#1;data_in = testData6[11388];
@(posedge clk);
#1;data_in = testData6[11389];
@(posedge clk);
#1;data_in = testData6[11390];
@(posedge clk);
#1;data_in = testData6[11391];
@(posedge clk);
#1;data_in = testData6[11392];
@(posedge clk);
#1;data_in = testData6[11393];
@(posedge clk);
#1;data_in = testData6[11394];
@(posedge clk);
#1;data_in = testData6[11395];
@(posedge clk);
#1;data_in = testData6[11396];
@(posedge clk);
#1;data_in = testData6[11397];
@(posedge clk);
#1;data_in = testData6[11398];
@(posedge clk);
#1;data_in = testData6[11399];
@(posedge clk);
#1;data_in = testData6[11400];
@(posedge clk);
#1;data_in = testData6[11401];
@(posedge clk);
#1;data_in = testData6[11402];
@(posedge clk);
#1;data_in = testData6[11403];
@(posedge clk);
#1;data_in = testData6[11404];
@(posedge clk);
#1;data_in = testData6[11405];
@(posedge clk);
#1;data_in = testData6[11406];
@(posedge clk);
#1;data_in = testData6[11407];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[11408]; 
@(posedge clk);
#1;data_in = testData6[11409];
@(posedge clk);
#1;data_in = testData6[11410];
@(posedge clk);
#1;data_in = testData6[11411];
@(posedge clk);
#1;data_in = testData6[11412];
@(posedge clk);
#1;data_in = testData6[11413];
@(posedge clk);
#1;data_in = testData6[11414];
@(posedge clk);
#1;data_in = testData6[11415];
@(posedge clk);
#1;data_in = testData6[11416];
@(posedge clk);
#1;data_in = testData6[11417];
@(posedge clk);
#1;data_in = testData6[11418];
@(posedge clk);
#1;data_in = testData6[11419];
@(posedge clk);
#1;data_in = testData6[11420];
@(posedge clk);
#1;data_in = testData6[11421];
@(posedge clk);
#1;data_in = testData6[11422];
@(posedge clk);
#1;data_in = testData6[11423];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[11424];
@(posedge clk);
#1;data_in = testData6[11425];
@(posedge clk);
#1;data_in = testData6[11426];
@(posedge clk);
#1;data_in = testData6[11427];
@(posedge clk);
#1;data_in = testData6[11428];
@(posedge clk);
#1;data_in = testData6[11429];
@(posedge clk);
#1;data_in = testData6[11430];
@(posedge clk);
#1;data_in = testData6[11431];
@(posedge clk);
#1;data_in = testData6[11432];
@(posedge clk);
#1;data_in = testData6[11433];
@(posedge clk);
#1;data_in = testData6[11434];
@(posedge clk);
#1;data_in = testData6[11435];
@(posedge clk);
#1;data_in = testData6[11436];
@(posedge clk);
#1;data_in = testData6[11437];
@(posedge clk);
#1;data_in = testData6[11438];
@(posedge clk);
#1;data_in = testData6[11439];
@(posedge clk);
#1;data_in = testData6[11440];
@(posedge clk);
#1;data_in = testData6[11441];
@(posedge clk);
#1;data_in = testData6[11442];
@(posedge clk);
#1;data_in = testData6[11443];
@(posedge clk);
#1;data_in = testData6[11444];
@(posedge clk);
#1;data_in = testData6[11445];
@(posedge clk);
#1;data_in = testData6[11446];
@(posedge clk);
#1;data_in = testData6[11447];
@(posedge clk);
#1;data_in = testData6[11448];
@(posedge clk);
#1;data_in = testData6[11449];
@(posedge clk);
#1;data_in = testData6[11450];
@(posedge clk);
#1;data_in = testData6[11451];
@(posedge clk);
#1;data_in = testData6[11452];
@(posedge clk);
#1;data_in = testData6[11453];
@(posedge clk);
#1;data_in = testData6[11454];
@(posedge clk);
#1;data_in = testData6[11455];
@(posedge clk);
#1;data_in = testData6[11456];
@(posedge clk);
#1;data_in = testData6[11457];
@(posedge clk);
#1;data_in = testData6[11458];
@(posedge clk);
#1;data_in = testData6[11459];
@(posedge clk);
#1;data_in = testData6[11460];
@(posedge clk);
#1;data_in = testData6[11461];
@(posedge clk);
#1;data_in = testData6[11462];
@(posedge clk);
#1;data_in = testData6[11463];
@(posedge clk);
#1;data_in = testData6[11464];
@(posedge clk);
#1;data_in = testData6[11465];
@(posedge clk);
#1;data_in = testData6[11466];
@(posedge clk);
#1;data_in = testData6[11467];
@(posedge clk);
#1;data_in = testData6[11468];
@(posedge clk);
#1;data_in = testData6[11469];
@(posedge clk);
#1;data_in = testData6[11470];
@(posedge clk);
#1;data_in = testData6[11471];
@(posedge clk);
#1;data_in = testData6[11472];
@(posedge clk);
#1;data_in = testData6[11473];
@(posedge clk);
#1;data_in = testData6[11474];
@(posedge clk);
#1;data_in = testData6[11475];
@(posedge clk);
#1;data_in = testData6[11476];
@(posedge clk);
#1;data_in = testData6[11477];
@(posedge clk);
#1;data_in = testData6[11478];
@(posedge clk);
#1;data_in = testData6[11479];
@(posedge clk);
#1;data_in = testData6[11480];
@(posedge clk);
#1;data_in = testData6[11481];
@(posedge clk);
#1;data_in = testData6[11482];
@(posedge clk);
#1;data_in = testData6[11483];
@(posedge clk);
#1;data_in = testData6[11484];
@(posedge clk);
#1;data_in = testData6[11485];
@(posedge clk);
#1;data_in = testData6[11486];
@(posedge clk);
#1;data_in = testData6[11487];
@(posedge clk);
#1;data_in = testData6[11488];
@(posedge clk);
#1;data_in = testData6[11489];
@(posedge clk);
#1;data_in = testData6[11490];
@(posedge clk);
#1;data_in = testData6[11491];
@(posedge clk);
#1;data_in = testData6[11492];
@(posedge clk);
#1;data_in = testData6[11493];
@(posedge clk);
#1;data_in = testData6[11494];
@(posedge clk);
#1;data_in = testData6[11495];
@(posedge clk);
#1;data_in = testData6[11496];
@(posedge clk);
#1;data_in = testData6[11497];
@(posedge clk);
#1;data_in = testData6[11498];
@(posedge clk);
#1;data_in = testData6[11499];
@(posedge clk);
#1;data_in = testData6[11500];
@(posedge clk);
#1;data_in = testData6[11501];
@(posedge clk);
#1;data_in = testData6[11502];
@(posedge clk);
#1;data_in = testData6[11503];
@(posedge clk);
#1;data_in = testData6[11504];
@(posedge clk);
#1;data_in = testData6[11505];
@(posedge clk);
#1;data_in = testData6[11506];
@(posedge clk);
#1;data_in = testData6[11507];
@(posedge clk);
#1;data_in = testData6[11508];
@(posedge clk);
#1;data_in = testData6[11509];
@(posedge clk);
#1;data_in = testData6[11510];
@(posedge clk);
#1;data_in = testData6[11511];
@(posedge clk);
#1;data_in = testData6[11512];
@(posedge clk);
#1;data_in = testData6[11513];
@(posedge clk);
#1;data_in = testData6[11514];
@(posedge clk);
#1;data_in = testData6[11515];
@(posedge clk);
#1;data_in = testData6[11516];
@(posedge clk);
#1;data_in = testData6[11517];
@(posedge clk);
#1;data_in = testData6[11518];
@(posedge clk);
#1;data_in = testData6[11519];
@(posedge clk);
#1;data_in = testData6[11520];
@(posedge clk);
#1;data_in = testData6[11521];
@(posedge clk);
#1;data_in = testData6[11522];
@(posedge clk);
#1;data_in = testData6[11523];
@(posedge clk);
#1;data_in = testData6[11524];
@(posedge clk);
#1;data_in = testData6[11525];
@(posedge clk);
#1;data_in = testData6[11526];
@(posedge clk);
#1;data_in = testData6[11527];
@(posedge clk);
#1;data_in = testData6[11528];
@(posedge clk);
#1;data_in = testData6[11529];
@(posedge clk);
#1;data_in = testData6[11530];
@(posedge clk);
#1;data_in = testData6[11531];
@(posedge clk);
#1;data_in = testData6[11532];
@(posedge clk);
#1;data_in = testData6[11533];
@(posedge clk);
#1;data_in = testData6[11534];
@(posedge clk);
#1;data_in = testData6[11535];
@(posedge clk);
#1;data_in = testData6[11536];
@(posedge clk);
#1;data_in = testData6[11537];
@(posedge clk);
#1;data_in = testData6[11538];
@(posedge clk);
#1;data_in = testData6[11539];
@(posedge clk);
#1;data_in = testData6[11540];
@(posedge clk);
#1;data_in = testData6[11541];
@(posedge clk);
#1;data_in = testData6[11542];
@(posedge clk);
#1;data_in = testData6[11543];
@(posedge clk);
#1;data_in = testData6[11544];
@(posedge clk);
#1;data_in = testData6[11545];
@(posedge clk);
#1;data_in = testData6[11546];
@(posedge clk);
#1;data_in = testData6[11547];
@(posedge clk);
#1;data_in = testData6[11548];
@(posedge clk);
#1;data_in = testData6[11549];
@(posedge clk);
#1;data_in = testData6[11550];
@(posedge clk);
#1;data_in = testData6[11551];
@(posedge clk);
#1;data_in = testData6[11552];
@(posedge clk);
#1;data_in = testData6[11553];
@(posedge clk);
#1;data_in = testData6[11554];
@(posedge clk);
#1;data_in = testData6[11555];
@(posedge clk);
#1;data_in = testData6[11556];
@(posedge clk);
#1;data_in = testData6[11557];
@(posedge clk);
#1;data_in = testData6[11558];
@(posedge clk);
#1;data_in = testData6[11559];
@(posedge clk);
#1;data_in = testData6[11560];
@(posedge clk);
#1;data_in = testData6[11561];
@(posedge clk);
#1;data_in = testData6[11562];
@(posedge clk);
#1;data_in = testData6[11563];
@(posedge clk);
#1;data_in = testData6[11564];
@(posedge clk);
#1;data_in = testData6[11565];
@(posedge clk);
#1;data_in = testData6[11566];
@(posedge clk);
#1;data_in = testData6[11567];
@(posedge clk);
#1;data_in = testData6[11568];
@(posedge clk);
#1;data_in = testData6[11569];
@(posedge clk);
#1;data_in = testData6[11570];
@(posedge clk);
#1;data_in = testData6[11571];
@(posedge clk);
#1;data_in = testData6[11572];
@(posedge clk);
#1;data_in = testData6[11573];
@(posedge clk);
#1;data_in = testData6[11574];
@(posedge clk);
#1;data_in = testData6[11575];
@(posedge clk);
#1;data_in = testData6[11576];
@(posedge clk);
#1;data_in = testData6[11577];
@(posedge clk);
#1;data_in = testData6[11578];
@(posedge clk);
#1;data_in = testData6[11579];
@(posedge clk);
#1;data_in = testData6[11580];
@(posedge clk);
#1;data_in = testData6[11581];
@(posedge clk);
#1;data_in = testData6[11582];
@(posedge clk);
#1;data_in = testData6[11583];
@(posedge clk);
#1;data_in = testData6[11584];
@(posedge clk);
#1;data_in = testData6[11585];
@(posedge clk);
#1;data_in = testData6[11586];
@(posedge clk);
#1;data_in = testData6[11587];
@(posedge clk);
#1;data_in = testData6[11588];
@(posedge clk);
#1;data_in = testData6[11589];
@(posedge clk);
#1;data_in = testData6[11590];
@(posedge clk);
#1;data_in = testData6[11591];
@(posedge clk);
#1;data_in = testData6[11592];
@(posedge clk);
#1;data_in = testData6[11593];
@(posedge clk);
#1;data_in = testData6[11594];
@(posedge clk);
#1;data_in = testData6[11595];
@(posedge clk);
#1;data_in = testData6[11596];
@(posedge clk);
#1;data_in = testData6[11597];
@(posedge clk);
#1;data_in = testData6[11598];
@(posedge clk);
#1;data_in = testData6[11599];
@(posedge clk);
#1;data_in = testData6[11600];
@(posedge clk);
#1;data_in = testData6[11601];
@(posedge clk);
#1;data_in = testData6[11602];
@(posedge clk);
#1;data_in = testData6[11603];
@(posedge clk);
#1;data_in = testData6[11604];
@(posedge clk);
#1;data_in = testData6[11605];
@(posedge clk);
#1;data_in = testData6[11606];
@(posedge clk);
#1;data_in = testData6[11607];
@(posedge clk);
#1;data_in = testData6[11608];
@(posedge clk);
#1;data_in = testData6[11609];
@(posedge clk);
#1;data_in = testData6[11610];
@(posedge clk);
#1;data_in = testData6[11611];
@(posedge clk);
#1;data_in = testData6[11612];
@(posedge clk);
#1;data_in = testData6[11613];
@(posedge clk);
#1;data_in = testData6[11614];
@(posedge clk);
#1;data_in = testData6[11615];
@(posedge clk);
#1;data_in = testData6[11616];
@(posedge clk);
#1;data_in = testData6[11617];
@(posedge clk);
#1;data_in = testData6[11618];
@(posedge clk);
#1;data_in = testData6[11619];
@(posedge clk);
#1;data_in = testData6[11620];
@(posedge clk);
#1;data_in = testData6[11621];
@(posedge clk);
#1;data_in = testData6[11622];
@(posedge clk);
#1;data_in = testData6[11623];
@(posedge clk);
#1;data_in = testData6[11624];
@(posedge clk);
#1;data_in = testData6[11625];
@(posedge clk);
#1;data_in = testData6[11626];
@(posedge clk);
#1;data_in = testData6[11627];
@(posedge clk);
#1;data_in = testData6[11628];
@(posedge clk);
#1;data_in = testData6[11629];
@(posedge clk);
#1;data_in = testData6[11630];
@(posedge clk);
#1;data_in = testData6[11631];
@(posedge clk);
#1;data_in = testData6[11632];
@(posedge clk);
#1;data_in = testData6[11633];
@(posedge clk);
#1;data_in = testData6[11634];
@(posedge clk);
#1;data_in = testData6[11635];
@(posedge clk);
#1;data_in = testData6[11636];
@(posedge clk);
#1;data_in = testData6[11637];
@(posedge clk);
#1;data_in = testData6[11638];
@(posedge clk);
#1;data_in = testData6[11639];
@(posedge clk);
#1;data_in = testData6[11640];
@(posedge clk);
#1;data_in = testData6[11641];
@(posedge clk);
#1;data_in = testData6[11642];
@(posedge clk);
#1;data_in = testData6[11643];
@(posedge clk);
#1;data_in = testData6[11644];
@(posedge clk);
#1;data_in = testData6[11645];
@(posedge clk);
#1;data_in = testData6[11646];
@(posedge clk);
#1;data_in = testData6[11647];
@(posedge clk);
#1;data_in = testData6[11648];
@(posedge clk);
#1;data_in = testData6[11649];
@(posedge clk);
#1;data_in = testData6[11650];
@(posedge clk);
#1;data_in = testData6[11651];
@(posedge clk);
#1;data_in = testData6[11652];
@(posedge clk);
#1;data_in = testData6[11653];
@(posedge clk);
#1;data_in = testData6[11654];
@(posedge clk);
#1;data_in = testData6[11655];
@(posedge clk);
#1;data_in = testData6[11656];
@(posedge clk);
#1;data_in = testData6[11657];
@(posedge clk);
#1;data_in = testData6[11658];
@(posedge clk);
#1;data_in = testData6[11659];
@(posedge clk);
#1;data_in = testData6[11660];
@(posedge clk);
#1;data_in = testData6[11661];
@(posedge clk);
#1;data_in = testData6[11662];
@(posedge clk);
#1;data_in = testData6[11663];
@(posedge clk);
#1;data_in = testData6[11664];
@(posedge clk);
#1;data_in = testData6[11665];
@(posedge clk);
#1;data_in = testData6[11666];
@(posedge clk);
#1;data_in = testData6[11667];
@(posedge clk);
#1;data_in = testData6[11668];
@(posedge clk);
#1;data_in = testData6[11669];
@(posedge clk);
#1;data_in = testData6[11670];
@(posedge clk);
#1;data_in = testData6[11671];
@(posedge clk);
#1;data_in = testData6[11672];
@(posedge clk);
#1;data_in = testData6[11673];
@(posedge clk);
#1;data_in = testData6[11674];
@(posedge clk);
#1;data_in = testData6[11675];
@(posedge clk);
#1;data_in = testData6[11676];
@(posedge clk);
#1;data_in = testData6[11677];
@(posedge clk);
#1;data_in = testData6[11678];
@(posedge clk);
#1;data_in = testData6[11679];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[11680]; 
@(posedge clk);
#1;data_in = testData6[11681];
@(posedge clk);
#1;data_in = testData6[11682];
@(posedge clk);
#1;data_in = testData6[11683];
@(posedge clk);
#1;data_in = testData6[11684];
@(posedge clk);
#1;data_in = testData6[11685];
@(posedge clk);
#1;data_in = testData6[11686];
@(posedge clk);
#1;data_in = testData6[11687];
@(posedge clk);
#1;data_in = testData6[11688];
@(posedge clk);
#1;data_in = testData6[11689];
@(posedge clk);
#1;data_in = testData6[11690];
@(posedge clk);
#1;data_in = testData6[11691];
@(posedge clk);
#1;data_in = testData6[11692];
@(posedge clk);
#1;data_in = testData6[11693];
@(posedge clk);
#1;data_in = testData6[11694];
@(posedge clk);
#1;data_in = testData6[11695];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[11696];
@(posedge clk);
#1;data_in = testData6[11697];
@(posedge clk);
#1;data_in = testData6[11698];
@(posedge clk);
#1;data_in = testData6[11699];
@(posedge clk);
#1;data_in = testData6[11700];
@(posedge clk);
#1;data_in = testData6[11701];
@(posedge clk);
#1;data_in = testData6[11702];
@(posedge clk);
#1;data_in = testData6[11703];
@(posedge clk);
#1;data_in = testData6[11704];
@(posedge clk);
#1;data_in = testData6[11705];
@(posedge clk);
#1;data_in = testData6[11706];
@(posedge clk);
#1;data_in = testData6[11707];
@(posedge clk);
#1;data_in = testData6[11708];
@(posedge clk);
#1;data_in = testData6[11709];
@(posedge clk);
#1;data_in = testData6[11710];
@(posedge clk);
#1;data_in = testData6[11711];
@(posedge clk);
#1;data_in = testData6[11712];
@(posedge clk);
#1;data_in = testData6[11713];
@(posedge clk);
#1;data_in = testData6[11714];
@(posedge clk);
#1;data_in = testData6[11715];
@(posedge clk);
#1;data_in = testData6[11716];
@(posedge clk);
#1;data_in = testData6[11717];
@(posedge clk);
#1;data_in = testData6[11718];
@(posedge clk);
#1;data_in = testData6[11719];
@(posedge clk);
#1;data_in = testData6[11720];
@(posedge clk);
#1;data_in = testData6[11721];
@(posedge clk);
#1;data_in = testData6[11722];
@(posedge clk);
#1;data_in = testData6[11723];
@(posedge clk);
#1;data_in = testData6[11724];
@(posedge clk);
#1;data_in = testData6[11725];
@(posedge clk);
#1;data_in = testData6[11726];
@(posedge clk);
#1;data_in = testData6[11727];
@(posedge clk);
#1;data_in = testData6[11728];
@(posedge clk);
#1;data_in = testData6[11729];
@(posedge clk);
#1;data_in = testData6[11730];
@(posedge clk);
#1;data_in = testData6[11731];
@(posedge clk);
#1;data_in = testData6[11732];
@(posedge clk);
#1;data_in = testData6[11733];
@(posedge clk);
#1;data_in = testData6[11734];
@(posedge clk);
#1;data_in = testData6[11735];
@(posedge clk);
#1;data_in = testData6[11736];
@(posedge clk);
#1;data_in = testData6[11737];
@(posedge clk);
#1;data_in = testData6[11738];
@(posedge clk);
#1;data_in = testData6[11739];
@(posedge clk);
#1;data_in = testData6[11740];
@(posedge clk);
#1;data_in = testData6[11741];
@(posedge clk);
#1;data_in = testData6[11742];
@(posedge clk);
#1;data_in = testData6[11743];
@(posedge clk);
#1;data_in = testData6[11744];
@(posedge clk);
#1;data_in = testData6[11745];
@(posedge clk);
#1;data_in = testData6[11746];
@(posedge clk);
#1;data_in = testData6[11747];
@(posedge clk);
#1;data_in = testData6[11748];
@(posedge clk);
#1;data_in = testData6[11749];
@(posedge clk);
#1;data_in = testData6[11750];
@(posedge clk);
#1;data_in = testData6[11751];
@(posedge clk);
#1;data_in = testData6[11752];
@(posedge clk);
#1;data_in = testData6[11753];
@(posedge clk);
#1;data_in = testData6[11754];
@(posedge clk);
#1;data_in = testData6[11755];
@(posedge clk);
#1;data_in = testData6[11756];
@(posedge clk);
#1;data_in = testData6[11757];
@(posedge clk);
#1;data_in = testData6[11758];
@(posedge clk);
#1;data_in = testData6[11759];
@(posedge clk);
#1;data_in = testData6[11760];
@(posedge clk);
#1;data_in = testData6[11761];
@(posedge clk);
#1;data_in = testData6[11762];
@(posedge clk);
#1;data_in = testData6[11763];
@(posedge clk);
#1;data_in = testData6[11764];
@(posedge clk);
#1;data_in = testData6[11765];
@(posedge clk);
#1;data_in = testData6[11766];
@(posedge clk);
#1;data_in = testData6[11767];
@(posedge clk);
#1;data_in = testData6[11768];
@(posedge clk);
#1;data_in = testData6[11769];
@(posedge clk);
#1;data_in = testData6[11770];
@(posedge clk);
#1;data_in = testData6[11771];
@(posedge clk);
#1;data_in = testData6[11772];
@(posedge clk);
#1;data_in = testData6[11773];
@(posedge clk);
#1;data_in = testData6[11774];
@(posedge clk);
#1;data_in = testData6[11775];
@(posedge clk);
#1;data_in = testData6[11776];
@(posedge clk);
#1;data_in = testData6[11777];
@(posedge clk);
#1;data_in = testData6[11778];
@(posedge clk);
#1;data_in = testData6[11779];
@(posedge clk);
#1;data_in = testData6[11780];
@(posedge clk);
#1;data_in = testData6[11781];
@(posedge clk);
#1;data_in = testData6[11782];
@(posedge clk);
#1;data_in = testData6[11783];
@(posedge clk);
#1;data_in = testData6[11784];
@(posedge clk);
#1;data_in = testData6[11785];
@(posedge clk);
#1;data_in = testData6[11786];
@(posedge clk);
#1;data_in = testData6[11787];
@(posedge clk);
#1;data_in = testData6[11788];
@(posedge clk);
#1;data_in = testData6[11789];
@(posedge clk);
#1;data_in = testData6[11790];
@(posedge clk);
#1;data_in = testData6[11791];
@(posedge clk);
#1;data_in = testData6[11792];
@(posedge clk);
#1;data_in = testData6[11793];
@(posedge clk);
#1;data_in = testData6[11794];
@(posedge clk);
#1;data_in = testData6[11795];
@(posedge clk);
#1;data_in = testData6[11796];
@(posedge clk);
#1;data_in = testData6[11797];
@(posedge clk);
#1;data_in = testData6[11798];
@(posedge clk);
#1;data_in = testData6[11799];
@(posedge clk);
#1;data_in = testData6[11800];
@(posedge clk);
#1;data_in = testData6[11801];
@(posedge clk);
#1;data_in = testData6[11802];
@(posedge clk);
#1;data_in = testData6[11803];
@(posedge clk);
#1;data_in = testData6[11804];
@(posedge clk);
#1;data_in = testData6[11805];
@(posedge clk);
#1;data_in = testData6[11806];
@(posedge clk);
#1;data_in = testData6[11807];
@(posedge clk);
#1;data_in = testData6[11808];
@(posedge clk);
#1;data_in = testData6[11809];
@(posedge clk);
#1;data_in = testData6[11810];
@(posedge clk);
#1;data_in = testData6[11811];
@(posedge clk);
#1;data_in = testData6[11812];
@(posedge clk);
#1;data_in = testData6[11813];
@(posedge clk);
#1;data_in = testData6[11814];
@(posedge clk);
#1;data_in = testData6[11815];
@(posedge clk);
#1;data_in = testData6[11816];
@(posedge clk);
#1;data_in = testData6[11817];
@(posedge clk);
#1;data_in = testData6[11818];
@(posedge clk);
#1;data_in = testData6[11819];
@(posedge clk);
#1;data_in = testData6[11820];
@(posedge clk);
#1;data_in = testData6[11821];
@(posedge clk);
#1;data_in = testData6[11822];
@(posedge clk);
#1;data_in = testData6[11823];
@(posedge clk);
#1;data_in = testData6[11824];
@(posedge clk);
#1;data_in = testData6[11825];
@(posedge clk);
#1;data_in = testData6[11826];
@(posedge clk);
#1;data_in = testData6[11827];
@(posedge clk);
#1;data_in = testData6[11828];
@(posedge clk);
#1;data_in = testData6[11829];
@(posedge clk);
#1;data_in = testData6[11830];
@(posedge clk);
#1;data_in = testData6[11831];
@(posedge clk);
#1;data_in = testData6[11832];
@(posedge clk);
#1;data_in = testData6[11833];
@(posedge clk);
#1;data_in = testData6[11834];
@(posedge clk);
#1;data_in = testData6[11835];
@(posedge clk);
#1;data_in = testData6[11836];
@(posedge clk);
#1;data_in = testData6[11837];
@(posedge clk);
#1;data_in = testData6[11838];
@(posedge clk);
#1;data_in = testData6[11839];
@(posedge clk);
#1;data_in = testData6[11840];
@(posedge clk);
#1;data_in = testData6[11841];
@(posedge clk);
#1;data_in = testData6[11842];
@(posedge clk);
#1;data_in = testData6[11843];
@(posedge clk);
#1;data_in = testData6[11844];
@(posedge clk);
#1;data_in = testData6[11845];
@(posedge clk);
#1;data_in = testData6[11846];
@(posedge clk);
#1;data_in = testData6[11847];
@(posedge clk);
#1;data_in = testData6[11848];
@(posedge clk);
#1;data_in = testData6[11849];
@(posedge clk);
#1;data_in = testData6[11850];
@(posedge clk);
#1;data_in = testData6[11851];
@(posedge clk);
#1;data_in = testData6[11852];
@(posedge clk);
#1;data_in = testData6[11853];
@(posedge clk);
#1;data_in = testData6[11854];
@(posedge clk);
#1;data_in = testData6[11855];
@(posedge clk);
#1;data_in = testData6[11856];
@(posedge clk);
#1;data_in = testData6[11857];
@(posedge clk);
#1;data_in = testData6[11858];
@(posedge clk);
#1;data_in = testData6[11859];
@(posedge clk);
#1;data_in = testData6[11860];
@(posedge clk);
#1;data_in = testData6[11861];
@(posedge clk);
#1;data_in = testData6[11862];
@(posedge clk);
#1;data_in = testData6[11863];
@(posedge clk);
#1;data_in = testData6[11864];
@(posedge clk);
#1;data_in = testData6[11865];
@(posedge clk);
#1;data_in = testData6[11866];
@(posedge clk);
#1;data_in = testData6[11867];
@(posedge clk);
#1;data_in = testData6[11868];
@(posedge clk);
#1;data_in = testData6[11869];
@(posedge clk);
#1;data_in = testData6[11870];
@(posedge clk);
#1;data_in = testData6[11871];
@(posedge clk);
#1;data_in = testData6[11872];
@(posedge clk);
#1;data_in = testData6[11873];
@(posedge clk);
#1;data_in = testData6[11874];
@(posedge clk);
#1;data_in = testData6[11875];
@(posedge clk);
#1;data_in = testData6[11876];
@(posedge clk);
#1;data_in = testData6[11877];
@(posedge clk);
#1;data_in = testData6[11878];
@(posedge clk);
#1;data_in = testData6[11879];
@(posedge clk);
#1;data_in = testData6[11880];
@(posedge clk);
#1;data_in = testData6[11881];
@(posedge clk);
#1;data_in = testData6[11882];
@(posedge clk);
#1;data_in = testData6[11883];
@(posedge clk);
#1;data_in = testData6[11884];
@(posedge clk);
#1;data_in = testData6[11885];
@(posedge clk);
#1;data_in = testData6[11886];
@(posedge clk);
#1;data_in = testData6[11887];
@(posedge clk);
#1;data_in = testData6[11888];
@(posedge clk);
#1;data_in = testData6[11889];
@(posedge clk);
#1;data_in = testData6[11890];
@(posedge clk);
#1;data_in = testData6[11891];
@(posedge clk);
#1;data_in = testData6[11892];
@(posedge clk);
#1;data_in = testData6[11893];
@(posedge clk);
#1;data_in = testData6[11894];
@(posedge clk);
#1;data_in = testData6[11895];
@(posedge clk);
#1;data_in = testData6[11896];
@(posedge clk);
#1;data_in = testData6[11897];
@(posedge clk);
#1;data_in = testData6[11898];
@(posedge clk);
#1;data_in = testData6[11899];
@(posedge clk);
#1;data_in = testData6[11900];
@(posedge clk);
#1;data_in = testData6[11901];
@(posedge clk);
#1;data_in = testData6[11902];
@(posedge clk);
#1;data_in = testData6[11903];
@(posedge clk);
#1;data_in = testData6[11904];
@(posedge clk);
#1;data_in = testData6[11905];
@(posedge clk);
#1;data_in = testData6[11906];
@(posedge clk);
#1;data_in = testData6[11907];
@(posedge clk);
#1;data_in = testData6[11908];
@(posedge clk);
#1;data_in = testData6[11909];
@(posedge clk);
#1;data_in = testData6[11910];
@(posedge clk);
#1;data_in = testData6[11911];
@(posedge clk);
#1;data_in = testData6[11912];
@(posedge clk);
#1;data_in = testData6[11913];
@(posedge clk);
#1;data_in = testData6[11914];
@(posedge clk);
#1;data_in = testData6[11915];
@(posedge clk);
#1;data_in = testData6[11916];
@(posedge clk);
#1;data_in = testData6[11917];
@(posedge clk);
#1;data_in = testData6[11918];
@(posedge clk);
#1;data_in = testData6[11919];
@(posedge clk);
#1;data_in = testData6[11920];
@(posedge clk);
#1;data_in = testData6[11921];
@(posedge clk);
#1;data_in = testData6[11922];
@(posedge clk);
#1;data_in = testData6[11923];
@(posedge clk);
#1;data_in = testData6[11924];
@(posedge clk);
#1;data_in = testData6[11925];
@(posedge clk);
#1;data_in = testData6[11926];
@(posedge clk);
#1;data_in = testData6[11927];
@(posedge clk);
#1;data_in = testData6[11928];
@(posedge clk);
#1;data_in = testData6[11929];
@(posedge clk);
#1;data_in = testData6[11930];
@(posedge clk);
#1;data_in = testData6[11931];
@(posedge clk);
#1;data_in = testData6[11932];
@(posedge clk);
#1;data_in = testData6[11933];
@(posedge clk);
#1;data_in = testData6[11934];
@(posedge clk);
#1;data_in = testData6[11935];
@(posedge clk);
#1;data_in = testData6[11936];
@(posedge clk);
#1;data_in = testData6[11937];
@(posedge clk);
#1;data_in = testData6[11938];
@(posedge clk);
#1;data_in = testData6[11939];
@(posedge clk);
#1;data_in = testData6[11940];
@(posedge clk);
#1;data_in = testData6[11941];
@(posedge clk);
#1;data_in = testData6[11942];
@(posedge clk);
#1;data_in = testData6[11943];
@(posedge clk);
#1;data_in = testData6[11944];
@(posedge clk);
#1;data_in = testData6[11945];
@(posedge clk);
#1;data_in = testData6[11946];
@(posedge clk);
#1;data_in = testData6[11947];
@(posedge clk);
#1;data_in = testData6[11948];
@(posedge clk);
#1;data_in = testData6[11949];
@(posedge clk);
#1;data_in = testData6[11950];
@(posedge clk);
#1;data_in = testData6[11951];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[11952]; 
@(posedge clk);
#1;data_in = testData6[11953];
@(posedge clk);
#1;data_in = testData6[11954];
@(posedge clk);
#1;data_in = testData6[11955];
@(posedge clk);
#1;data_in = testData6[11956];
@(posedge clk);
#1;data_in = testData6[11957];
@(posedge clk);
#1;data_in = testData6[11958];
@(posedge clk);
#1;data_in = testData6[11959];
@(posedge clk);
#1;data_in = testData6[11960];
@(posedge clk);
#1;data_in = testData6[11961];
@(posedge clk);
#1;data_in = testData6[11962];
@(posedge clk);
#1;data_in = testData6[11963];
@(posedge clk);
#1;data_in = testData6[11964];
@(posedge clk);
#1;data_in = testData6[11965];
@(posedge clk);
#1;data_in = testData6[11966];
@(posedge clk);
#1;data_in = testData6[11967];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[11968];
@(posedge clk);
#1;data_in = testData6[11969];
@(posedge clk);
#1;data_in = testData6[11970];
@(posedge clk);
#1;data_in = testData6[11971];
@(posedge clk);
#1;data_in = testData6[11972];
@(posedge clk);
#1;data_in = testData6[11973];
@(posedge clk);
#1;data_in = testData6[11974];
@(posedge clk);
#1;data_in = testData6[11975];
@(posedge clk);
#1;data_in = testData6[11976];
@(posedge clk);
#1;data_in = testData6[11977];
@(posedge clk);
#1;data_in = testData6[11978];
@(posedge clk);
#1;data_in = testData6[11979];
@(posedge clk);
#1;data_in = testData6[11980];
@(posedge clk);
#1;data_in = testData6[11981];
@(posedge clk);
#1;data_in = testData6[11982];
@(posedge clk);
#1;data_in = testData6[11983];
@(posedge clk);
#1;data_in = testData6[11984];
@(posedge clk);
#1;data_in = testData6[11985];
@(posedge clk);
#1;data_in = testData6[11986];
@(posedge clk);
#1;data_in = testData6[11987];
@(posedge clk);
#1;data_in = testData6[11988];
@(posedge clk);
#1;data_in = testData6[11989];
@(posedge clk);
#1;data_in = testData6[11990];
@(posedge clk);
#1;data_in = testData6[11991];
@(posedge clk);
#1;data_in = testData6[11992];
@(posedge clk);
#1;data_in = testData6[11993];
@(posedge clk);
#1;data_in = testData6[11994];
@(posedge clk);
#1;data_in = testData6[11995];
@(posedge clk);
#1;data_in = testData6[11996];
@(posedge clk);
#1;data_in = testData6[11997];
@(posedge clk);
#1;data_in = testData6[11998];
@(posedge clk);
#1;data_in = testData6[11999];
@(posedge clk);
#1;data_in = testData6[12000];
@(posedge clk);
#1;data_in = testData6[12001];
@(posedge clk);
#1;data_in = testData6[12002];
@(posedge clk);
#1;data_in = testData6[12003];
@(posedge clk);
#1;data_in = testData6[12004];
@(posedge clk);
#1;data_in = testData6[12005];
@(posedge clk);
#1;data_in = testData6[12006];
@(posedge clk);
#1;data_in = testData6[12007];
@(posedge clk);
#1;data_in = testData6[12008];
@(posedge clk);
#1;data_in = testData6[12009];
@(posedge clk);
#1;data_in = testData6[12010];
@(posedge clk);
#1;data_in = testData6[12011];
@(posedge clk);
#1;data_in = testData6[12012];
@(posedge clk);
#1;data_in = testData6[12013];
@(posedge clk);
#1;data_in = testData6[12014];
@(posedge clk);
#1;data_in = testData6[12015];
@(posedge clk);
#1;data_in = testData6[12016];
@(posedge clk);
#1;data_in = testData6[12017];
@(posedge clk);
#1;data_in = testData6[12018];
@(posedge clk);
#1;data_in = testData6[12019];
@(posedge clk);
#1;data_in = testData6[12020];
@(posedge clk);
#1;data_in = testData6[12021];
@(posedge clk);
#1;data_in = testData6[12022];
@(posedge clk);
#1;data_in = testData6[12023];
@(posedge clk);
#1;data_in = testData6[12024];
@(posedge clk);
#1;data_in = testData6[12025];
@(posedge clk);
#1;data_in = testData6[12026];
@(posedge clk);
#1;data_in = testData6[12027];
@(posedge clk);
#1;data_in = testData6[12028];
@(posedge clk);
#1;data_in = testData6[12029];
@(posedge clk);
#1;data_in = testData6[12030];
@(posedge clk);
#1;data_in = testData6[12031];
@(posedge clk);
#1;data_in = testData6[12032];
@(posedge clk);
#1;data_in = testData6[12033];
@(posedge clk);
#1;data_in = testData6[12034];
@(posedge clk);
#1;data_in = testData6[12035];
@(posedge clk);
#1;data_in = testData6[12036];
@(posedge clk);
#1;data_in = testData6[12037];
@(posedge clk);
#1;data_in = testData6[12038];
@(posedge clk);
#1;data_in = testData6[12039];
@(posedge clk);
#1;data_in = testData6[12040];
@(posedge clk);
#1;data_in = testData6[12041];
@(posedge clk);
#1;data_in = testData6[12042];
@(posedge clk);
#1;data_in = testData6[12043];
@(posedge clk);
#1;data_in = testData6[12044];
@(posedge clk);
#1;data_in = testData6[12045];
@(posedge clk);
#1;data_in = testData6[12046];
@(posedge clk);
#1;data_in = testData6[12047];
@(posedge clk);
#1;data_in = testData6[12048];
@(posedge clk);
#1;data_in = testData6[12049];
@(posedge clk);
#1;data_in = testData6[12050];
@(posedge clk);
#1;data_in = testData6[12051];
@(posedge clk);
#1;data_in = testData6[12052];
@(posedge clk);
#1;data_in = testData6[12053];
@(posedge clk);
#1;data_in = testData6[12054];
@(posedge clk);
#1;data_in = testData6[12055];
@(posedge clk);
#1;data_in = testData6[12056];
@(posedge clk);
#1;data_in = testData6[12057];
@(posedge clk);
#1;data_in = testData6[12058];
@(posedge clk);
#1;data_in = testData6[12059];
@(posedge clk);
#1;data_in = testData6[12060];
@(posedge clk);
#1;data_in = testData6[12061];
@(posedge clk);
#1;data_in = testData6[12062];
@(posedge clk);
#1;data_in = testData6[12063];
@(posedge clk);
#1;data_in = testData6[12064];
@(posedge clk);
#1;data_in = testData6[12065];
@(posedge clk);
#1;data_in = testData6[12066];
@(posedge clk);
#1;data_in = testData6[12067];
@(posedge clk);
#1;data_in = testData6[12068];
@(posedge clk);
#1;data_in = testData6[12069];
@(posedge clk);
#1;data_in = testData6[12070];
@(posedge clk);
#1;data_in = testData6[12071];
@(posedge clk);
#1;data_in = testData6[12072];
@(posedge clk);
#1;data_in = testData6[12073];
@(posedge clk);
#1;data_in = testData6[12074];
@(posedge clk);
#1;data_in = testData6[12075];
@(posedge clk);
#1;data_in = testData6[12076];
@(posedge clk);
#1;data_in = testData6[12077];
@(posedge clk);
#1;data_in = testData6[12078];
@(posedge clk);
#1;data_in = testData6[12079];
@(posedge clk);
#1;data_in = testData6[12080];
@(posedge clk);
#1;data_in = testData6[12081];
@(posedge clk);
#1;data_in = testData6[12082];
@(posedge clk);
#1;data_in = testData6[12083];
@(posedge clk);
#1;data_in = testData6[12084];
@(posedge clk);
#1;data_in = testData6[12085];
@(posedge clk);
#1;data_in = testData6[12086];
@(posedge clk);
#1;data_in = testData6[12087];
@(posedge clk);
#1;data_in = testData6[12088];
@(posedge clk);
#1;data_in = testData6[12089];
@(posedge clk);
#1;data_in = testData6[12090];
@(posedge clk);
#1;data_in = testData6[12091];
@(posedge clk);
#1;data_in = testData6[12092];
@(posedge clk);
#1;data_in = testData6[12093];
@(posedge clk);
#1;data_in = testData6[12094];
@(posedge clk);
#1;data_in = testData6[12095];
@(posedge clk);
#1;data_in = testData6[12096];
@(posedge clk);
#1;data_in = testData6[12097];
@(posedge clk);
#1;data_in = testData6[12098];
@(posedge clk);
#1;data_in = testData6[12099];
@(posedge clk);
#1;data_in = testData6[12100];
@(posedge clk);
#1;data_in = testData6[12101];
@(posedge clk);
#1;data_in = testData6[12102];
@(posedge clk);
#1;data_in = testData6[12103];
@(posedge clk);
#1;data_in = testData6[12104];
@(posedge clk);
#1;data_in = testData6[12105];
@(posedge clk);
#1;data_in = testData6[12106];
@(posedge clk);
#1;data_in = testData6[12107];
@(posedge clk);
#1;data_in = testData6[12108];
@(posedge clk);
#1;data_in = testData6[12109];
@(posedge clk);
#1;data_in = testData6[12110];
@(posedge clk);
#1;data_in = testData6[12111];
@(posedge clk);
#1;data_in = testData6[12112];
@(posedge clk);
#1;data_in = testData6[12113];
@(posedge clk);
#1;data_in = testData6[12114];
@(posedge clk);
#1;data_in = testData6[12115];
@(posedge clk);
#1;data_in = testData6[12116];
@(posedge clk);
#1;data_in = testData6[12117];
@(posedge clk);
#1;data_in = testData6[12118];
@(posedge clk);
#1;data_in = testData6[12119];
@(posedge clk);
#1;data_in = testData6[12120];
@(posedge clk);
#1;data_in = testData6[12121];
@(posedge clk);
#1;data_in = testData6[12122];
@(posedge clk);
#1;data_in = testData6[12123];
@(posedge clk);
#1;data_in = testData6[12124];
@(posedge clk);
#1;data_in = testData6[12125];
@(posedge clk);
#1;data_in = testData6[12126];
@(posedge clk);
#1;data_in = testData6[12127];
@(posedge clk);
#1;data_in = testData6[12128];
@(posedge clk);
#1;data_in = testData6[12129];
@(posedge clk);
#1;data_in = testData6[12130];
@(posedge clk);
#1;data_in = testData6[12131];
@(posedge clk);
#1;data_in = testData6[12132];
@(posedge clk);
#1;data_in = testData6[12133];
@(posedge clk);
#1;data_in = testData6[12134];
@(posedge clk);
#1;data_in = testData6[12135];
@(posedge clk);
#1;data_in = testData6[12136];
@(posedge clk);
#1;data_in = testData6[12137];
@(posedge clk);
#1;data_in = testData6[12138];
@(posedge clk);
#1;data_in = testData6[12139];
@(posedge clk);
#1;data_in = testData6[12140];
@(posedge clk);
#1;data_in = testData6[12141];
@(posedge clk);
#1;data_in = testData6[12142];
@(posedge clk);
#1;data_in = testData6[12143];
@(posedge clk);
#1;data_in = testData6[12144];
@(posedge clk);
#1;data_in = testData6[12145];
@(posedge clk);
#1;data_in = testData6[12146];
@(posedge clk);
#1;data_in = testData6[12147];
@(posedge clk);
#1;data_in = testData6[12148];
@(posedge clk);
#1;data_in = testData6[12149];
@(posedge clk);
#1;data_in = testData6[12150];
@(posedge clk);
#1;data_in = testData6[12151];
@(posedge clk);
#1;data_in = testData6[12152];
@(posedge clk);
#1;data_in = testData6[12153];
@(posedge clk);
#1;data_in = testData6[12154];
@(posedge clk);
#1;data_in = testData6[12155];
@(posedge clk);
#1;data_in = testData6[12156];
@(posedge clk);
#1;data_in = testData6[12157];
@(posedge clk);
#1;data_in = testData6[12158];
@(posedge clk);
#1;data_in = testData6[12159];
@(posedge clk);
#1;data_in = testData6[12160];
@(posedge clk);
#1;data_in = testData6[12161];
@(posedge clk);
#1;data_in = testData6[12162];
@(posedge clk);
#1;data_in = testData6[12163];
@(posedge clk);
#1;data_in = testData6[12164];
@(posedge clk);
#1;data_in = testData6[12165];
@(posedge clk);
#1;data_in = testData6[12166];
@(posedge clk);
#1;data_in = testData6[12167];
@(posedge clk);
#1;data_in = testData6[12168];
@(posedge clk);
#1;data_in = testData6[12169];
@(posedge clk);
#1;data_in = testData6[12170];
@(posedge clk);
#1;data_in = testData6[12171];
@(posedge clk);
#1;data_in = testData6[12172];
@(posedge clk);
#1;data_in = testData6[12173];
@(posedge clk);
#1;data_in = testData6[12174];
@(posedge clk);
#1;data_in = testData6[12175];
@(posedge clk);
#1;data_in = testData6[12176];
@(posedge clk);
#1;data_in = testData6[12177];
@(posedge clk);
#1;data_in = testData6[12178];
@(posedge clk);
#1;data_in = testData6[12179];
@(posedge clk);
#1;data_in = testData6[12180];
@(posedge clk);
#1;data_in = testData6[12181];
@(posedge clk);
#1;data_in = testData6[12182];
@(posedge clk);
#1;data_in = testData6[12183];
@(posedge clk);
#1;data_in = testData6[12184];
@(posedge clk);
#1;data_in = testData6[12185];
@(posedge clk);
#1;data_in = testData6[12186];
@(posedge clk);
#1;data_in = testData6[12187];
@(posedge clk);
#1;data_in = testData6[12188];
@(posedge clk);
#1;data_in = testData6[12189];
@(posedge clk);
#1;data_in = testData6[12190];
@(posedge clk);
#1;data_in = testData6[12191];
@(posedge clk);
#1;data_in = testData6[12192];
@(posedge clk);
#1;data_in = testData6[12193];
@(posedge clk);
#1;data_in = testData6[12194];
@(posedge clk);
#1;data_in = testData6[12195];
@(posedge clk);
#1;data_in = testData6[12196];
@(posedge clk);
#1;data_in = testData6[12197];
@(posedge clk);
#1;data_in = testData6[12198];
@(posedge clk);
#1;data_in = testData6[12199];
@(posedge clk);
#1;data_in = testData6[12200];
@(posedge clk);
#1;data_in = testData6[12201];
@(posedge clk);
#1;data_in = testData6[12202];
@(posedge clk);
#1;data_in = testData6[12203];
@(posedge clk);
#1;data_in = testData6[12204];
@(posedge clk);
#1;data_in = testData6[12205];
@(posedge clk);
#1;data_in = testData6[12206];
@(posedge clk);
#1;data_in = testData6[12207];
@(posedge clk);
#1;data_in = testData6[12208];
@(posedge clk);
#1;data_in = testData6[12209];
@(posedge clk);
#1;data_in = testData6[12210];
@(posedge clk);
#1;data_in = testData6[12211];
@(posedge clk);
#1;data_in = testData6[12212];
@(posedge clk);
#1;data_in = testData6[12213];
@(posedge clk);
#1;data_in = testData6[12214];
@(posedge clk);
#1;data_in = testData6[12215];
@(posedge clk);
#1;data_in = testData6[12216];
@(posedge clk);
#1;data_in = testData6[12217];
@(posedge clk);
#1;data_in = testData6[12218];
@(posedge clk);
#1;data_in = testData6[12219];
@(posedge clk);
#1;data_in = testData6[12220];
@(posedge clk);
#1;data_in = testData6[12221];
@(posedge clk);
#1;data_in = testData6[12222];
@(posedge clk);
#1;data_in = testData6[12223];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[12224]; 
@(posedge clk);
#1;data_in = testData6[12225];
@(posedge clk);
#1;data_in = testData6[12226];
@(posedge clk);
#1;data_in = testData6[12227];
@(posedge clk);
#1;data_in = testData6[12228];
@(posedge clk);
#1;data_in = testData6[12229];
@(posedge clk);
#1;data_in = testData6[12230];
@(posedge clk);
#1;data_in = testData6[12231];
@(posedge clk);
#1;data_in = testData6[12232];
@(posedge clk);
#1;data_in = testData6[12233];
@(posedge clk);
#1;data_in = testData6[12234];
@(posedge clk);
#1;data_in = testData6[12235];
@(posedge clk);
#1;data_in = testData6[12236];
@(posedge clk);
#1;data_in = testData6[12237];
@(posedge clk);
#1;data_in = testData6[12238];
@(posedge clk);
#1;data_in = testData6[12239];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[12240];
@(posedge clk);
#1;data_in = testData6[12241];
@(posedge clk);
#1;data_in = testData6[12242];
@(posedge clk);
#1;data_in = testData6[12243];
@(posedge clk);
#1;data_in = testData6[12244];
@(posedge clk);
#1;data_in = testData6[12245];
@(posedge clk);
#1;data_in = testData6[12246];
@(posedge clk);
#1;data_in = testData6[12247];
@(posedge clk);
#1;data_in = testData6[12248];
@(posedge clk);
#1;data_in = testData6[12249];
@(posedge clk);
#1;data_in = testData6[12250];
@(posedge clk);
#1;data_in = testData6[12251];
@(posedge clk);
#1;data_in = testData6[12252];
@(posedge clk);
#1;data_in = testData6[12253];
@(posedge clk);
#1;data_in = testData6[12254];
@(posedge clk);
#1;data_in = testData6[12255];
@(posedge clk);
#1;data_in = testData6[12256];
@(posedge clk);
#1;data_in = testData6[12257];
@(posedge clk);
#1;data_in = testData6[12258];
@(posedge clk);
#1;data_in = testData6[12259];
@(posedge clk);
#1;data_in = testData6[12260];
@(posedge clk);
#1;data_in = testData6[12261];
@(posedge clk);
#1;data_in = testData6[12262];
@(posedge clk);
#1;data_in = testData6[12263];
@(posedge clk);
#1;data_in = testData6[12264];
@(posedge clk);
#1;data_in = testData6[12265];
@(posedge clk);
#1;data_in = testData6[12266];
@(posedge clk);
#1;data_in = testData6[12267];
@(posedge clk);
#1;data_in = testData6[12268];
@(posedge clk);
#1;data_in = testData6[12269];
@(posedge clk);
#1;data_in = testData6[12270];
@(posedge clk);
#1;data_in = testData6[12271];
@(posedge clk);
#1;data_in = testData6[12272];
@(posedge clk);
#1;data_in = testData6[12273];
@(posedge clk);
#1;data_in = testData6[12274];
@(posedge clk);
#1;data_in = testData6[12275];
@(posedge clk);
#1;data_in = testData6[12276];
@(posedge clk);
#1;data_in = testData6[12277];
@(posedge clk);
#1;data_in = testData6[12278];
@(posedge clk);
#1;data_in = testData6[12279];
@(posedge clk);
#1;data_in = testData6[12280];
@(posedge clk);
#1;data_in = testData6[12281];
@(posedge clk);
#1;data_in = testData6[12282];
@(posedge clk);
#1;data_in = testData6[12283];
@(posedge clk);
#1;data_in = testData6[12284];
@(posedge clk);
#1;data_in = testData6[12285];
@(posedge clk);
#1;data_in = testData6[12286];
@(posedge clk);
#1;data_in = testData6[12287];
@(posedge clk);
#1;data_in = testData6[12288];
@(posedge clk);
#1;data_in = testData6[12289];
@(posedge clk);
#1;data_in = testData6[12290];
@(posedge clk);
#1;data_in = testData6[12291];
@(posedge clk);
#1;data_in = testData6[12292];
@(posedge clk);
#1;data_in = testData6[12293];
@(posedge clk);
#1;data_in = testData6[12294];
@(posedge clk);
#1;data_in = testData6[12295];
@(posedge clk);
#1;data_in = testData6[12296];
@(posedge clk);
#1;data_in = testData6[12297];
@(posedge clk);
#1;data_in = testData6[12298];
@(posedge clk);
#1;data_in = testData6[12299];
@(posedge clk);
#1;data_in = testData6[12300];
@(posedge clk);
#1;data_in = testData6[12301];
@(posedge clk);
#1;data_in = testData6[12302];
@(posedge clk);
#1;data_in = testData6[12303];
@(posedge clk);
#1;data_in = testData6[12304];
@(posedge clk);
#1;data_in = testData6[12305];
@(posedge clk);
#1;data_in = testData6[12306];
@(posedge clk);
#1;data_in = testData6[12307];
@(posedge clk);
#1;data_in = testData6[12308];
@(posedge clk);
#1;data_in = testData6[12309];
@(posedge clk);
#1;data_in = testData6[12310];
@(posedge clk);
#1;data_in = testData6[12311];
@(posedge clk);
#1;data_in = testData6[12312];
@(posedge clk);
#1;data_in = testData6[12313];
@(posedge clk);
#1;data_in = testData6[12314];
@(posedge clk);
#1;data_in = testData6[12315];
@(posedge clk);
#1;data_in = testData6[12316];
@(posedge clk);
#1;data_in = testData6[12317];
@(posedge clk);
#1;data_in = testData6[12318];
@(posedge clk);
#1;data_in = testData6[12319];
@(posedge clk);
#1;data_in = testData6[12320];
@(posedge clk);
#1;data_in = testData6[12321];
@(posedge clk);
#1;data_in = testData6[12322];
@(posedge clk);
#1;data_in = testData6[12323];
@(posedge clk);
#1;data_in = testData6[12324];
@(posedge clk);
#1;data_in = testData6[12325];
@(posedge clk);
#1;data_in = testData6[12326];
@(posedge clk);
#1;data_in = testData6[12327];
@(posedge clk);
#1;data_in = testData6[12328];
@(posedge clk);
#1;data_in = testData6[12329];
@(posedge clk);
#1;data_in = testData6[12330];
@(posedge clk);
#1;data_in = testData6[12331];
@(posedge clk);
#1;data_in = testData6[12332];
@(posedge clk);
#1;data_in = testData6[12333];
@(posedge clk);
#1;data_in = testData6[12334];
@(posedge clk);
#1;data_in = testData6[12335];
@(posedge clk);
#1;data_in = testData6[12336];
@(posedge clk);
#1;data_in = testData6[12337];
@(posedge clk);
#1;data_in = testData6[12338];
@(posedge clk);
#1;data_in = testData6[12339];
@(posedge clk);
#1;data_in = testData6[12340];
@(posedge clk);
#1;data_in = testData6[12341];
@(posedge clk);
#1;data_in = testData6[12342];
@(posedge clk);
#1;data_in = testData6[12343];
@(posedge clk);
#1;data_in = testData6[12344];
@(posedge clk);
#1;data_in = testData6[12345];
@(posedge clk);
#1;data_in = testData6[12346];
@(posedge clk);
#1;data_in = testData6[12347];
@(posedge clk);
#1;data_in = testData6[12348];
@(posedge clk);
#1;data_in = testData6[12349];
@(posedge clk);
#1;data_in = testData6[12350];
@(posedge clk);
#1;data_in = testData6[12351];
@(posedge clk);
#1;data_in = testData6[12352];
@(posedge clk);
#1;data_in = testData6[12353];
@(posedge clk);
#1;data_in = testData6[12354];
@(posedge clk);
#1;data_in = testData6[12355];
@(posedge clk);
#1;data_in = testData6[12356];
@(posedge clk);
#1;data_in = testData6[12357];
@(posedge clk);
#1;data_in = testData6[12358];
@(posedge clk);
#1;data_in = testData6[12359];
@(posedge clk);
#1;data_in = testData6[12360];
@(posedge clk);
#1;data_in = testData6[12361];
@(posedge clk);
#1;data_in = testData6[12362];
@(posedge clk);
#1;data_in = testData6[12363];
@(posedge clk);
#1;data_in = testData6[12364];
@(posedge clk);
#1;data_in = testData6[12365];
@(posedge clk);
#1;data_in = testData6[12366];
@(posedge clk);
#1;data_in = testData6[12367];
@(posedge clk);
#1;data_in = testData6[12368];
@(posedge clk);
#1;data_in = testData6[12369];
@(posedge clk);
#1;data_in = testData6[12370];
@(posedge clk);
#1;data_in = testData6[12371];
@(posedge clk);
#1;data_in = testData6[12372];
@(posedge clk);
#1;data_in = testData6[12373];
@(posedge clk);
#1;data_in = testData6[12374];
@(posedge clk);
#1;data_in = testData6[12375];
@(posedge clk);
#1;data_in = testData6[12376];
@(posedge clk);
#1;data_in = testData6[12377];
@(posedge clk);
#1;data_in = testData6[12378];
@(posedge clk);
#1;data_in = testData6[12379];
@(posedge clk);
#1;data_in = testData6[12380];
@(posedge clk);
#1;data_in = testData6[12381];
@(posedge clk);
#1;data_in = testData6[12382];
@(posedge clk);
#1;data_in = testData6[12383];
@(posedge clk);
#1;data_in = testData6[12384];
@(posedge clk);
#1;data_in = testData6[12385];
@(posedge clk);
#1;data_in = testData6[12386];
@(posedge clk);
#1;data_in = testData6[12387];
@(posedge clk);
#1;data_in = testData6[12388];
@(posedge clk);
#1;data_in = testData6[12389];
@(posedge clk);
#1;data_in = testData6[12390];
@(posedge clk);
#1;data_in = testData6[12391];
@(posedge clk);
#1;data_in = testData6[12392];
@(posedge clk);
#1;data_in = testData6[12393];
@(posedge clk);
#1;data_in = testData6[12394];
@(posedge clk);
#1;data_in = testData6[12395];
@(posedge clk);
#1;data_in = testData6[12396];
@(posedge clk);
#1;data_in = testData6[12397];
@(posedge clk);
#1;data_in = testData6[12398];
@(posedge clk);
#1;data_in = testData6[12399];
@(posedge clk);
#1;data_in = testData6[12400];
@(posedge clk);
#1;data_in = testData6[12401];
@(posedge clk);
#1;data_in = testData6[12402];
@(posedge clk);
#1;data_in = testData6[12403];
@(posedge clk);
#1;data_in = testData6[12404];
@(posedge clk);
#1;data_in = testData6[12405];
@(posedge clk);
#1;data_in = testData6[12406];
@(posedge clk);
#1;data_in = testData6[12407];
@(posedge clk);
#1;data_in = testData6[12408];
@(posedge clk);
#1;data_in = testData6[12409];
@(posedge clk);
#1;data_in = testData6[12410];
@(posedge clk);
#1;data_in = testData6[12411];
@(posedge clk);
#1;data_in = testData6[12412];
@(posedge clk);
#1;data_in = testData6[12413];
@(posedge clk);
#1;data_in = testData6[12414];
@(posedge clk);
#1;data_in = testData6[12415];
@(posedge clk);
#1;data_in = testData6[12416];
@(posedge clk);
#1;data_in = testData6[12417];
@(posedge clk);
#1;data_in = testData6[12418];
@(posedge clk);
#1;data_in = testData6[12419];
@(posedge clk);
#1;data_in = testData6[12420];
@(posedge clk);
#1;data_in = testData6[12421];
@(posedge clk);
#1;data_in = testData6[12422];
@(posedge clk);
#1;data_in = testData6[12423];
@(posedge clk);
#1;data_in = testData6[12424];
@(posedge clk);
#1;data_in = testData6[12425];
@(posedge clk);
#1;data_in = testData6[12426];
@(posedge clk);
#1;data_in = testData6[12427];
@(posedge clk);
#1;data_in = testData6[12428];
@(posedge clk);
#1;data_in = testData6[12429];
@(posedge clk);
#1;data_in = testData6[12430];
@(posedge clk);
#1;data_in = testData6[12431];
@(posedge clk);
#1;data_in = testData6[12432];
@(posedge clk);
#1;data_in = testData6[12433];
@(posedge clk);
#1;data_in = testData6[12434];
@(posedge clk);
#1;data_in = testData6[12435];
@(posedge clk);
#1;data_in = testData6[12436];
@(posedge clk);
#1;data_in = testData6[12437];
@(posedge clk);
#1;data_in = testData6[12438];
@(posedge clk);
#1;data_in = testData6[12439];
@(posedge clk);
#1;data_in = testData6[12440];
@(posedge clk);
#1;data_in = testData6[12441];
@(posedge clk);
#1;data_in = testData6[12442];
@(posedge clk);
#1;data_in = testData6[12443];
@(posedge clk);
#1;data_in = testData6[12444];
@(posedge clk);
#1;data_in = testData6[12445];
@(posedge clk);
#1;data_in = testData6[12446];
@(posedge clk);
#1;data_in = testData6[12447];
@(posedge clk);
#1;data_in = testData6[12448];
@(posedge clk);
#1;data_in = testData6[12449];
@(posedge clk);
#1;data_in = testData6[12450];
@(posedge clk);
#1;data_in = testData6[12451];
@(posedge clk);
#1;data_in = testData6[12452];
@(posedge clk);
#1;data_in = testData6[12453];
@(posedge clk);
#1;data_in = testData6[12454];
@(posedge clk);
#1;data_in = testData6[12455];
@(posedge clk);
#1;data_in = testData6[12456];
@(posedge clk);
#1;data_in = testData6[12457];
@(posedge clk);
#1;data_in = testData6[12458];
@(posedge clk);
#1;data_in = testData6[12459];
@(posedge clk);
#1;data_in = testData6[12460];
@(posedge clk);
#1;data_in = testData6[12461];
@(posedge clk);
#1;data_in = testData6[12462];
@(posedge clk);
#1;data_in = testData6[12463];
@(posedge clk);
#1;data_in = testData6[12464];
@(posedge clk);
#1;data_in = testData6[12465];
@(posedge clk);
#1;data_in = testData6[12466];
@(posedge clk);
#1;data_in = testData6[12467];
@(posedge clk);
#1;data_in = testData6[12468];
@(posedge clk);
#1;data_in = testData6[12469];
@(posedge clk);
#1;data_in = testData6[12470];
@(posedge clk);
#1;data_in = testData6[12471];
@(posedge clk);
#1;data_in = testData6[12472];
@(posedge clk);
#1;data_in = testData6[12473];
@(posedge clk);
#1;data_in = testData6[12474];
@(posedge clk);
#1;data_in = testData6[12475];
@(posedge clk);
#1;data_in = testData6[12476];
@(posedge clk);
#1;data_in = testData6[12477];
@(posedge clk);
#1;data_in = testData6[12478];
@(posedge clk);
#1;data_in = testData6[12479];
@(posedge clk);
#1;data_in = testData6[12480];
@(posedge clk);
#1;data_in = testData6[12481];
@(posedge clk);
#1;data_in = testData6[12482];
@(posedge clk);
#1;data_in = testData6[12483];
@(posedge clk);
#1;data_in = testData6[12484];
@(posedge clk);
#1;data_in = testData6[12485];
@(posedge clk);
#1;data_in = testData6[12486];
@(posedge clk);
#1;data_in = testData6[12487];
@(posedge clk);
#1;data_in = testData6[12488];
@(posedge clk);
#1;data_in = testData6[12489];
@(posedge clk);
#1;data_in = testData6[12490];
@(posedge clk);
#1;data_in = testData6[12491];
@(posedge clk);
#1;data_in = testData6[12492];
@(posedge clk);
#1;data_in = testData6[12493];
@(posedge clk);
#1;data_in = testData6[12494];
@(posedge clk);
#1;data_in = testData6[12495];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[12496]; 
@(posedge clk);
#1;data_in = testData6[12497];
@(posedge clk);
#1;data_in = testData6[12498];
@(posedge clk);
#1;data_in = testData6[12499];
@(posedge clk);
#1;data_in = testData6[12500];
@(posedge clk);
#1;data_in = testData6[12501];
@(posedge clk);
#1;data_in = testData6[12502];
@(posedge clk);
#1;data_in = testData6[12503];
@(posedge clk);
#1;data_in = testData6[12504];
@(posedge clk);
#1;data_in = testData6[12505];
@(posedge clk);
#1;data_in = testData6[12506];
@(posedge clk);
#1;data_in = testData6[12507];
@(posedge clk);
#1;data_in = testData6[12508];
@(posedge clk);
#1;data_in = testData6[12509];
@(posedge clk);
#1;data_in = testData6[12510];
@(posedge clk);
#1;data_in = testData6[12511];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[12512];
@(posedge clk);
#1;data_in = testData6[12513];
@(posedge clk);
#1;data_in = testData6[12514];
@(posedge clk);
#1;data_in = testData6[12515];
@(posedge clk);
#1;data_in = testData6[12516];
@(posedge clk);
#1;data_in = testData6[12517];
@(posedge clk);
#1;data_in = testData6[12518];
@(posedge clk);
#1;data_in = testData6[12519];
@(posedge clk);
#1;data_in = testData6[12520];
@(posedge clk);
#1;data_in = testData6[12521];
@(posedge clk);
#1;data_in = testData6[12522];
@(posedge clk);
#1;data_in = testData6[12523];
@(posedge clk);
#1;data_in = testData6[12524];
@(posedge clk);
#1;data_in = testData6[12525];
@(posedge clk);
#1;data_in = testData6[12526];
@(posedge clk);
#1;data_in = testData6[12527];
@(posedge clk);
#1;data_in = testData6[12528];
@(posedge clk);
#1;data_in = testData6[12529];
@(posedge clk);
#1;data_in = testData6[12530];
@(posedge clk);
#1;data_in = testData6[12531];
@(posedge clk);
#1;data_in = testData6[12532];
@(posedge clk);
#1;data_in = testData6[12533];
@(posedge clk);
#1;data_in = testData6[12534];
@(posedge clk);
#1;data_in = testData6[12535];
@(posedge clk);
#1;data_in = testData6[12536];
@(posedge clk);
#1;data_in = testData6[12537];
@(posedge clk);
#1;data_in = testData6[12538];
@(posedge clk);
#1;data_in = testData6[12539];
@(posedge clk);
#1;data_in = testData6[12540];
@(posedge clk);
#1;data_in = testData6[12541];
@(posedge clk);
#1;data_in = testData6[12542];
@(posedge clk);
#1;data_in = testData6[12543];
@(posedge clk);
#1;data_in = testData6[12544];
@(posedge clk);
#1;data_in = testData6[12545];
@(posedge clk);
#1;data_in = testData6[12546];
@(posedge clk);
#1;data_in = testData6[12547];
@(posedge clk);
#1;data_in = testData6[12548];
@(posedge clk);
#1;data_in = testData6[12549];
@(posedge clk);
#1;data_in = testData6[12550];
@(posedge clk);
#1;data_in = testData6[12551];
@(posedge clk);
#1;data_in = testData6[12552];
@(posedge clk);
#1;data_in = testData6[12553];
@(posedge clk);
#1;data_in = testData6[12554];
@(posedge clk);
#1;data_in = testData6[12555];
@(posedge clk);
#1;data_in = testData6[12556];
@(posedge clk);
#1;data_in = testData6[12557];
@(posedge clk);
#1;data_in = testData6[12558];
@(posedge clk);
#1;data_in = testData6[12559];
@(posedge clk);
#1;data_in = testData6[12560];
@(posedge clk);
#1;data_in = testData6[12561];
@(posedge clk);
#1;data_in = testData6[12562];
@(posedge clk);
#1;data_in = testData6[12563];
@(posedge clk);
#1;data_in = testData6[12564];
@(posedge clk);
#1;data_in = testData6[12565];
@(posedge clk);
#1;data_in = testData6[12566];
@(posedge clk);
#1;data_in = testData6[12567];
@(posedge clk);
#1;data_in = testData6[12568];
@(posedge clk);
#1;data_in = testData6[12569];
@(posedge clk);
#1;data_in = testData6[12570];
@(posedge clk);
#1;data_in = testData6[12571];
@(posedge clk);
#1;data_in = testData6[12572];
@(posedge clk);
#1;data_in = testData6[12573];
@(posedge clk);
#1;data_in = testData6[12574];
@(posedge clk);
#1;data_in = testData6[12575];
@(posedge clk);
#1;data_in = testData6[12576];
@(posedge clk);
#1;data_in = testData6[12577];
@(posedge clk);
#1;data_in = testData6[12578];
@(posedge clk);
#1;data_in = testData6[12579];
@(posedge clk);
#1;data_in = testData6[12580];
@(posedge clk);
#1;data_in = testData6[12581];
@(posedge clk);
#1;data_in = testData6[12582];
@(posedge clk);
#1;data_in = testData6[12583];
@(posedge clk);
#1;data_in = testData6[12584];
@(posedge clk);
#1;data_in = testData6[12585];
@(posedge clk);
#1;data_in = testData6[12586];
@(posedge clk);
#1;data_in = testData6[12587];
@(posedge clk);
#1;data_in = testData6[12588];
@(posedge clk);
#1;data_in = testData6[12589];
@(posedge clk);
#1;data_in = testData6[12590];
@(posedge clk);
#1;data_in = testData6[12591];
@(posedge clk);
#1;data_in = testData6[12592];
@(posedge clk);
#1;data_in = testData6[12593];
@(posedge clk);
#1;data_in = testData6[12594];
@(posedge clk);
#1;data_in = testData6[12595];
@(posedge clk);
#1;data_in = testData6[12596];
@(posedge clk);
#1;data_in = testData6[12597];
@(posedge clk);
#1;data_in = testData6[12598];
@(posedge clk);
#1;data_in = testData6[12599];
@(posedge clk);
#1;data_in = testData6[12600];
@(posedge clk);
#1;data_in = testData6[12601];
@(posedge clk);
#1;data_in = testData6[12602];
@(posedge clk);
#1;data_in = testData6[12603];
@(posedge clk);
#1;data_in = testData6[12604];
@(posedge clk);
#1;data_in = testData6[12605];
@(posedge clk);
#1;data_in = testData6[12606];
@(posedge clk);
#1;data_in = testData6[12607];
@(posedge clk);
#1;data_in = testData6[12608];
@(posedge clk);
#1;data_in = testData6[12609];
@(posedge clk);
#1;data_in = testData6[12610];
@(posedge clk);
#1;data_in = testData6[12611];
@(posedge clk);
#1;data_in = testData6[12612];
@(posedge clk);
#1;data_in = testData6[12613];
@(posedge clk);
#1;data_in = testData6[12614];
@(posedge clk);
#1;data_in = testData6[12615];
@(posedge clk);
#1;data_in = testData6[12616];
@(posedge clk);
#1;data_in = testData6[12617];
@(posedge clk);
#1;data_in = testData6[12618];
@(posedge clk);
#1;data_in = testData6[12619];
@(posedge clk);
#1;data_in = testData6[12620];
@(posedge clk);
#1;data_in = testData6[12621];
@(posedge clk);
#1;data_in = testData6[12622];
@(posedge clk);
#1;data_in = testData6[12623];
@(posedge clk);
#1;data_in = testData6[12624];
@(posedge clk);
#1;data_in = testData6[12625];
@(posedge clk);
#1;data_in = testData6[12626];
@(posedge clk);
#1;data_in = testData6[12627];
@(posedge clk);
#1;data_in = testData6[12628];
@(posedge clk);
#1;data_in = testData6[12629];
@(posedge clk);
#1;data_in = testData6[12630];
@(posedge clk);
#1;data_in = testData6[12631];
@(posedge clk);
#1;data_in = testData6[12632];
@(posedge clk);
#1;data_in = testData6[12633];
@(posedge clk);
#1;data_in = testData6[12634];
@(posedge clk);
#1;data_in = testData6[12635];
@(posedge clk);
#1;data_in = testData6[12636];
@(posedge clk);
#1;data_in = testData6[12637];
@(posedge clk);
#1;data_in = testData6[12638];
@(posedge clk);
#1;data_in = testData6[12639];
@(posedge clk);
#1;data_in = testData6[12640];
@(posedge clk);
#1;data_in = testData6[12641];
@(posedge clk);
#1;data_in = testData6[12642];
@(posedge clk);
#1;data_in = testData6[12643];
@(posedge clk);
#1;data_in = testData6[12644];
@(posedge clk);
#1;data_in = testData6[12645];
@(posedge clk);
#1;data_in = testData6[12646];
@(posedge clk);
#1;data_in = testData6[12647];
@(posedge clk);
#1;data_in = testData6[12648];
@(posedge clk);
#1;data_in = testData6[12649];
@(posedge clk);
#1;data_in = testData6[12650];
@(posedge clk);
#1;data_in = testData6[12651];
@(posedge clk);
#1;data_in = testData6[12652];
@(posedge clk);
#1;data_in = testData6[12653];
@(posedge clk);
#1;data_in = testData6[12654];
@(posedge clk);
#1;data_in = testData6[12655];
@(posedge clk);
#1;data_in = testData6[12656];
@(posedge clk);
#1;data_in = testData6[12657];
@(posedge clk);
#1;data_in = testData6[12658];
@(posedge clk);
#1;data_in = testData6[12659];
@(posedge clk);
#1;data_in = testData6[12660];
@(posedge clk);
#1;data_in = testData6[12661];
@(posedge clk);
#1;data_in = testData6[12662];
@(posedge clk);
#1;data_in = testData6[12663];
@(posedge clk);
#1;data_in = testData6[12664];
@(posedge clk);
#1;data_in = testData6[12665];
@(posedge clk);
#1;data_in = testData6[12666];
@(posedge clk);
#1;data_in = testData6[12667];
@(posedge clk);
#1;data_in = testData6[12668];
@(posedge clk);
#1;data_in = testData6[12669];
@(posedge clk);
#1;data_in = testData6[12670];
@(posedge clk);
#1;data_in = testData6[12671];
@(posedge clk);
#1;data_in = testData6[12672];
@(posedge clk);
#1;data_in = testData6[12673];
@(posedge clk);
#1;data_in = testData6[12674];
@(posedge clk);
#1;data_in = testData6[12675];
@(posedge clk);
#1;data_in = testData6[12676];
@(posedge clk);
#1;data_in = testData6[12677];
@(posedge clk);
#1;data_in = testData6[12678];
@(posedge clk);
#1;data_in = testData6[12679];
@(posedge clk);
#1;data_in = testData6[12680];
@(posedge clk);
#1;data_in = testData6[12681];
@(posedge clk);
#1;data_in = testData6[12682];
@(posedge clk);
#1;data_in = testData6[12683];
@(posedge clk);
#1;data_in = testData6[12684];
@(posedge clk);
#1;data_in = testData6[12685];
@(posedge clk);
#1;data_in = testData6[12686];
@(posedge clk);
#1;data_in = testData6[12687];
@(posedge clk);
#1;data_in = testData6[12688];
@(posedge clk);
#1;data_in = testData6[12689];
@(posedge clk);
#1;data_in = testData6[12690];
@(posedge clk);
#1;data_in = testData6[12691];
@(posedge clk);
#1;data_in = testData6[12692];
@(posedge clk);
#1;data_in = testData6[12693];
@(posedge clk);
#1;data_in = testData6[12694];
@(posedge clk);
#1;data_in = testData6[12695];
@(posedge clk);
#1;data_in = testData6[12696];
@(posedge clk);
#1;data_in = testData6[12697];
@(posedge clk);
#1;data_in = testData6[12698];
@(posedge clk);
#1;data_in = testData6[12699];
@(posedge clk);
#1;data_in = testData6[12700];
@(posedge clk);
#1;data_in = testData6[12701];
@(posedge clk);
#1;data_in = testData6[12702];
@(posedge clk);
#1;data_in = testData6[12703];
@(posedge clk);
#1;data_in = testData6[12704];
@(posedge clk);
#1;data_in = testData6[12705];
@(posedge clk);
#1;data_in = testData6[12706];
@(posedge clk);
#1;data_in = testData6[12707];
@(posedge clk);
#1;data_in = testData6[12708];
@(posedge clk);
#1;data_in = testData6[12709];
@(posedge clk);
#1;data_in = testData6[12710];
@(posedge clk);
#1;data_in = testData6[12711];
@(posedge clk);
#1;data_in = testData6[12712];
@(posedge clk);
#1;data_in = testData6[12713];
@(posedge clk);
#1;data_in = testData6[12714];
@(posedge clk);
#1;data_in = testData6[12715];
@(posedge clk);
#1;data_in = testData6[12716];
@(posedge clk);
#1;data_in = testData6[12717];
@(posedge clk);
#1;data_in = testData6[12718];
@(posedge clk);
#1;data_in = testData6[12719];
@(posedge clk);
#1;data_in = testData6[12720];
@(posedge clk);
#1;data_in = testData6[12721];
@(posedge clk);
#1;data_in = testData6[12722];
@(posedge clk);
#1;data_in = testData6[12723];
@(posedge clk);
#1;data_in = testData6[12724];
@(posedge clk);
#1;data_in = testData6[12725];
@(posedge clk);
#1;data_in = testData6[12726];
@(posedge clk);
#1;data_in = testData6[12727];
@(posedge clk);
#1;data_in = testData6[12728];
@(posedge clk);
#1;data_in = testData6[12729];
@(posedge clk);
#1;data_in = testData6[12730];
@(posedge clk);
#1;data_in = testData6[12731];
@(posedge clk);
#1;data_in = testData6[12732];
@(posedge clk);
#1;data_in = testData6[12733];
@(posedge clk);
#1;data_in = testData6[12734];
@(posedge clk);
#1;data_in = testData6[12735];
@(posedge clk);
#1;data_in = testData6[12736];
@(posedge clk);
#1;data_in = testData6[12737];
@(posedge clk);
#1;data_in = testData6[12738];
@(posedge clk);
#1;data_in = testData6[12739];
@(posedge clk);
#1;data_in = testData6[12740];
@(posedge clk);
#1;data_in = testData6[12741];
@(posedge clk);
#1;data_in = testData6[12742];
@(posedge clk);
#1;data_in = testData6[12743];
@(posedge clk);
#1;data_in = testData6[12744];
@(posedge clk);
#1;data_in = testData6[12745];
@(posedge clk);
#1;data_in = testData6[12746];
@(posedge clk);
#1;data_in = testData6[12747];
@(posedge clk);
#1;data_in = testData6[12748];
@(posedge clk);
#1;data_in = testData6[12749];
@(posedge clk);
#1;data_in = testData6[12750];
@(posedge clk);
#1;data_in = testData6[12751];
@(posedge clk);
#1;data_in = testData6[12752];
@(posedge clk);
#1;data_in = testData6[12753];
@(posedge clk);
#1;data_in = testData6[12754];
@(posedge clk);
#1;data_in = testData6[12755];
@(posedge clk);
#1;data_in = testData6[12756];
@(posedge clk);
#1;data_in = testData6[12757];
@(posedge clk);
#1;data_in = testData6[12758];
@(posedge clk);
#1;data_in = testData6[12759];
@(posedge clk);
#1;data_in = testData6[12760];
@(posedge clk);
#1;data_in = testData6[12761];
@(posedge clk);
#1;data_in = testData6[12762];
@(posedge clk);
#1;data_in = testData6[12763];
@(posedge clk);
#1;data_in = testData6[12764];
@(posedge clk);
#1;data_in = testData6[12765];
@(posedge clk);
#1;data_in = testData6[12766];
@(posedge clk);
#1;data_in = testData6[12767];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[12768]; 
@(posedge clk);
#1;data_in = testData6[12769];
@(posedge clk);
#1;data_in = testData6[12770];
@(posedge clk);
#1;data_in = testData6[12771];
@(posedge clk);
#1;data_in = testData6[12772];
@(posedge clk);
#1;data_in = testData6[12773];
@(posedge clk);
#1;data_in = testData6[12774];
@(posedge clk);
#1;data_in = testData6[12775];
@(posedge clk);
#1;data_in = testData6[12776];
@(posedge clk);
#1;data_in = testData6[12777];
@(posedge clk);
#1;data_in = testData6[12778];
@(posedge clk);
#1;data_in = testData6[12779];
@(posedge clk);
#1;data_in = testData6[12780];
@(posedge clk);
#1;data_in = testData6[12781];
@(posedge clk);
#1;data_in = testData6[12782];
@(posedge clk);
#1;data_in = testData6[12783];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[12784];
@(posedge clk);
#1;data_in = testData6[12785];
@(posedge clk);
#1;data_in = testData6[12786];
@(posedge clk);
#1;data_in = testData6[12787];
@(posedge clk);
#1;data_in = testData6[12788];
@(posedge clk);
#1;data_in = testData6[12789];
@(posedge clk);
#1;data_in = testData6[12790];
@(posedge clk);
#1;data_in = testData6[12791];
@(posedge clk);
#1;data_in = testData6[12792];
@(posedge clk);
#1;data_in = testData6[12793];
@(posedge clk);
#1;data_in = testData6[12794];
@(posedge clk);
#1;data_in = testData6[12795];
@(posedge clk);
#1;data_in = testData6[12796];
@(posedge clk);
#1;data_in = testData6[12797];
@(posedge clk);
#1;data_in = testData6[12798];
@(posedge clk);
#1;data_in = testData6[12799];
@(posedge clk);
#1;data_in = testData6[12800];
@(posedge clk);
#1;data_in = testData6[12801];
@(posedge clk);
#1;data_in = testData6[12802];
@(posedge clk);
#1;data_in = testData6[12803];
@(posedge clk);
#1;data_in = testData6[12804];
@(posedge clk);
#1;data_in = testData6[12805];
@(posedge clk);
#1;data_in = testData6[12806];
@(posedge clk);
#1;data_in = testData6[12807];
@(posedge clk);
#1;data_in = testData6[12808];
@(posedge clk);
#1;data_in = testData6[12809];
@(posedge clk);
#1;data_in = testData6[12810];
@(posedge clk);
#1;data_in = testData6[12811];
@(posedge clk);
#1;data_in = testData6[12812];
@(posedge clk);
#1;data_in = testData6[12813];
@(posedge clk);
#1;data_in = testData6[12814];
@(posedge clk);
#1;data_in = testData6[12815];
@(posedge clk);
#1;data_in = testData6[12816];
@(posedge clk);
#1;data_in = testData6[12817];
@(posedge clk);
#1;data_in = testData6[12818];
@(posedge clk);
#1;data_in = testData6[12819];
@(posedge clk);
#1;data_in = testData6[12820];
@(posedge clk);
#1;data_in = testData6[12821];
@(posedge clk);
#1;data_in = testData6[12822];
@(posedge clk);
#1;data_in = testData6[12823];
@(posedge clk);
#1;data_in = testData6[12824];
@(posedge clk);
#1;data_in = testData6[12825];
@(posedge clk);
#1;data_in = testData6[12826];
@(posedge clk);
#1;data_in = testData6[12827];
@(posedge clk);
#1;data_in = testData6[12828];
@(posedge clk);
#1;data_in = testData6[12829];
@(posedge clk);
#1;data_in = testData6[12830];
@(posedge clk);
#1;data_in = testData6[12831];
@(posedge clk);
#1;data_in = testData6[12832];
@(posedge clk);
#1;data_in = testData6[12833];
@(posedge clk);
#1;data_in = testData6[12834];
@(posedge clk);
#1;data_in = testData6[12835];
@(posedge clk);
#1;data_in = testData6[12836];
@(posedge clk);
#1;data_in = testData6[12837];
@(posedge clk);
#1;data_in = testData6[12838];
@(posedge clk);
#1;data_in = testData6[12839];
@(posedge clk);
#1;data_in = testData6[12840];
@(posedge clk);
#1;data_in = testData6[12841];
@(posedge clk);
#1;data_in = testData6[12842];
@(posedge clk);
#1;data_in = testData6[12843];
@(posedge clk);
#1;data_in = testData6[12844];
@(posedge clk);
#1;data_in = testData6[12845];
@(posedge clk);
#1;data_in = testData6[12846];
@(posedge clk);
#1;data_in = testData6[12847];
@(posedge clk);
#1;data_in = testData6[12848];
@(posedge clk);
#1;data_in = testData6[12849];
@(posedge clk);
#1;data_in = testData6[12850];
@(posedge clk);
#1;data_in = testData6[12851];
@(posedge clk);
#1;data_in = testData6[12852];
@(posedge clk);
#1;data_in = testData6[12853];
@(posedge clk);
#1;data_in = testData6[12854];
@(posedge clk);
#1;data_in = testData6[12855];
@(posedge clk);
#1;data_in = testData6[12856];
@(posedge clk);
#1;data_in = testData6[12857];
@(posedge clk);
#1;data_in = testData6[12858];
@(posedge clk);
#1;data_in = testData6[12859];
@(posedge clk);
#1;data_in = testData6[12860];
@(posedge clk);
#1;data_in = testData6[12861];
@(posedge clk);
#1;data_in = testData6[12862];
@(posedge clk);
#1;data_in = testData6[12863];
@(posedge clk);
#1;data_in = testData6[12864];
@(posedge clk);
#1;data_in = testData6[12865];
@(posedge clk);
#1;data_in = testData6[12866];
@(posedge clk);
#1;data_in = testData6[12867];
@(posedge clk);
#1;data_in = testData6[12868];
@(posedge clk);
#1;data_in = testData6[12869];
@(posedge clk);
#1;data_in = testData6[12870];
@(posedge clk);
#1;data_in = testData6[12871];
@(posedge clk);
#1;data_in = testData6[12872];
@(posedge clk);
#1;data_in = testData6[12873];
@(posedge clk);
#1;data_in = testData6[12874];
@(posedge clk);
#1;data_in = testData6[12875];
@(posedge clk);
#1;data_in = testData6[12876];
@(posedge clk);
#1;data_in = testData6[12877];
@(posedge clk);
#1;data_in = testData6[12878];
@(posedge clk);
#1;data_in = testData6[12879];
@(posedge clk);
#1;data_in = testData6[12880];
@(posedge clk);
#1;data_in = testData6[12881];
@(posedge clk);
#1;data_in = testData6[12882];
@(posedge clk);
#1;data_in = testData6[12883];
@(posedge clk);
#1;data_in = testData6[12884];
@(posedge clk);
#1;data_in = testData6[12885];
@(posedge clk);
#1;data_in = testData6[12886];
@(posedge clk);
#1;data_in = testData6[12887];
@(posedge clk);
#1;data_in = testData6[12888];
@(posedge clk);
#1;data_in = testData6[12889];
@(posedge clk);
#1;data_in = testData6[12890];
@(posedge clk);
#1;data_in = testData6[12891];
@(posedge clk);
#1;data_in = testData6[12892];
@(posedge clk);
#1;data_in = testData6[12893];
@(posedge clk);
#1;data_in = testData6[12894];
@(posedge clk);
#1;data_in = testData6[12895];
@(posedge clk);
#1;data_in = testData6[12896];
@(posedge clk);
#1;data_in = testData6[12897];
@(posedge clk);
#1;data_in = testData6[12898];
@(posedge clk);
#1;data_in = testData6[12899];
@(posedge clk);
#1;data_in = testData6[12900];
@(posedge clk);
#1;data_in = testData6[12901];
@(posedge clk);
#1;data_in = testData6[12902];
@(posedge clk);
#1;data_in = testData6[12903];
@(posedge clk);
#1;data_in = testData6[12904];
@(posedge clk);
#1;data_in = testData6[12905];
@(posedge clk);
#1;data_in = testData6[12906];
@(posedge clk);
#1;data_in = testData6[12907];
@(posedge clk);
#1;data_in = testData6[12908];
@(posedge clk);
#1;data_in = testData6[12909];
@(posedge clk);
#1;data_in = testData6[12910];
@(posedge clk);
#1;data_in = testData6[12911];
@(posedge clk);
#1;data_in = testData6[12912];
@(posedge clk);
#1;data_in = testData6[12913];
@(posedge clk);
#1;data_in = testData6[12914];
@(posedge clk);
#1;data_in = testData6[12915];
@(posedge clk);
#1;data_in = testData6[12916];
@(posedge clk);
#1;data_in = testData6[12917];
@(posedge clk);
#1;data_in = testData6[12918];
@(posedge clk);
#1;data_in = testData6[12919];
@(posedge clk);
#1;data_in = testData6[12920];
@(posedge clk);
#1;data_in = testData6[12921];
@(posedge clk);
#1;data_in = testData6[12922];
@(posedge clk);
#1;data_in = testData6[12923];
@(posedge clk);
#1;data_in = testData6[12924];
@(posedge clk);
#1;data_in = testData6[12925];
@(posedge clk);
#1;data_in = testData6[12926];
@(posedge clk);
#1;data_in = testData6[12927];
@(posedge clk);
#1;data_in = testData6[12928];
@(posedge clk);
#1;data_in = testData6[12929];
@(posedge clk);
#1;data_in = testData6[12930];
@(posedge clk);
#1;data_in = testData6[12931];
@(posedge clk);
#1;data_in = testData6[12932];
@(posedge clk);
#1;data_in = testData6[12933];
@(posedge clk);
#1;data_in = testData6[12934];
@(posedge clk);
#1;data_in = testData6[12935];
@(posedge clk);
#1;data_in = testData6[12936];
@(posedge clk);
#1;data_in = testData6[12937];
@(posedge clk);
#1;data_in = testData6[12938];
@(posedge clk);
#1;data_in = testData6[12939];
@(posedge clk);
#1;data_in = testData6[12940];
@(posedge clk);
#1;data_in = testData6[12941];
@(posedge clk);
#1;data_in = testData6[12942];
@(posedge clk);
#1;data_in = testData6[12943];
@(posedge clk);
#1;data_in = testData6[12944];
@(posedge clk);
#1;data_in = testData6[12945];
@(posedge clk);
#1;data_in = testData6[12946];
@(posedge clk);
#1;data_in = testData6[12947];
@(posedge clk);
#1;data_in = testData6[12948];
@(posedge clk);
#1;data_in = testData6[12949];
@(posedge clk);
#1;data_in = testData6[12950];
@(posedge clk);
#1;data_in = testData6[12951];
@(posedge clk);
#1;data_in = testData6[12952];
@(posedge clk);
#1;data_in = testData6[12953];
@(posedge clk);
#1;data_in = testData6[12954];
@(posedge clk);
#1;data_in = testData6[12955];
@(posedge clk);
#1;data_in = testData6[12956];
@(posedge clk);
#1;data_in = testData6[12957];
@(posedge clk);
#1;data_in = testData6[12958];
@(posedge clk);
#1;data_in = testData6[12959];
@(posedge clk);
#1;data_in = testData6[12960];
@(posedge clk);
#1;data_in = testData6[12961];
@(posedge clk);
#1;data_in = testData6[12962];
@(posedge clk);
#1;data_in = testData6[12963];
@(posedge clk);
#1;data_in = testData6[12964];
@(posedge clk);
#1;data_in = testData6[12965];
@(posedge clk);
#1;data_in = testData6[12966];
@(posedge clk);
#1;data_in = testData6[12967];
@(posedge clk);
#1;data_in = testData6[12968];
@(posedge clk);
#1;data_in = testData6[12969];
@(posedge clk);
#1;data_in = testData6[12970];
@(posedge clk);
#1;data_in = testData6[12971];
@(posedge clk);
#1;data_in = testData6[12972];
@(posedge clk);
#1;data_in = testData6[12973];
@(posedge clk);
#1;data_in = testData6[12974];
@(posedge clk);
#1;data_in = testData6[12975];
@(posedge clk);
#1;data_in = testData6[12976];
@(posedge clk);
#1;data_in = testData6[12977];
@(posedge clk);
#1;data_in = testData6[12978];
@(posedge clk);
#1;data_in = testData6[12979];
@(posedge clk);
#1;data_in = testData6[12980];
@(posedge clk);
#1;data_in = testData6[12981];
@(posedge clk);
#1;data_in = testData6[12982];
@(posedge clk);
#1;data_in = testData6[12983];
@(posedge clk);
#1;data_in = testData6[12984];
@(posedge clk);
#1;data_in = testData6[12985];
@(posedge clk);
#1;data_in = testData6[12986];
@(posedge clk);
#1;data_in = testData6[12987];
@(posedge clk);
#1;data_in = testData6[12988];
@(posedge clk);
#1;data_in = testData6[12989];
@(posedge clk);
#1;data_in = testData6[12990];
@(posedge clk);
#1;data_in = testData6[12991];
@(posedge clk);
#1;data_in = testData6[12992];
@(posedge clk);
#1;data_in = testData6[12993];
@(posedge clk);
#1;data_in = testData6[12994];
@(posedge clk);
#1;data_in = testData6[12995];
@(posedge clk);
#1;data_in = testData6[12996];
@(posedge clk);
#1;data_in = testData6[12997];
@(posedge clk);
#1;data_in = testData6[12998];
@(posedge clk);
#1;data_in = testData6[12999];
@(posedge clk);
#1;data_in = testData6[13000];
@(posedge clk);
#1;data_in = testData6[13001];
@(posedge clk);
#1;data_in = testData6[13002];
@(posedge clk);
#1;data_in = testData6[13003];
@(posedge clk);
#1;data_in = testData6[13004];
@(posedge clk);
#1;data_in = testData6[13005];
@(posedge clk);
#1;data_in = testData6[13006];
@(posedge clk);
#1;data_in = testData6[13007];
@(posedge clk);
#1;data_in = testData6[13008];
@(posedge clk);
#1;data_in = testData6[13009];
@(posedge clk);
#1;data_in = testData6[13010];
@(posedge clk);
#1;data_in = testData6[13011];
@(posedge clk);
#1;data_in = testData6[13012];
@(posedge clk);
#1;data_in = testData6[13013];
@(posedge clk);
#1;data_in = testData6[13014];
@(posedge clk);
#1;data_in = testData6[13015];
@(posedge clk);
#1;data_in = testData6[13016];
@(posedge clk);
#1;data_in = testData6[13017];
@(posedge clk);
#1;data_in = testData6[13018];
@(posedge clk);
#1;data_in = testData6[13019];
@(posedge clk);
#1;data_in = testData6[13020];
@(posedge clk);
#1;data_in = testData6[13021];
@(posedge clk);
#1;data_in = testData6[13022];
@(posedge clk);
#1;data_in = testData6[13023];
@(posedge clk);
#1;data_in = testData6[13024];
@(posedge clk);
#1;data_in = testData6[13025];
@(posedge clk);
#1;data_in = testData6[13026];
@(posedge clk);
#1;data_in = testData6[13027];
@(posedge clk);
#1;data_in = testData6[13028];
@(posedge clk);
#1;data_in = testData6[13029];
@(posedge clk);
#1;data_in = testData6[13030];
@(posedge clk);
#1;data_in = testData6[13031];
@(posedge clk);
#1;data_in = testData6[13032];
@(posedge clk);
#1;data_in = testData6[13033];
@(posedge clk);
#1;data_in = testData6[13034];
@(posedge clk);
#1;data_in = testData6[13035];
@(posedge clk);
#1;data_in = testData6[13036];
@(posedge clk);
#1;data_in = testData6[13037];
@(posedge clk);
#1;data_in = testData6[13038];
@(posedge clk);
#1;data_in = testData6[13039];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[13040]; 
@(posedge clk);
#1;data_in = testData6[13041];
@(posedge clk);
#1;data_in = testData6[13042];
@(posedge clk);
#1;data_in = testData6[13043];
@(posedge clk);
#1;data_in = testData6[13044];
@(posedge clk);
#1;data_in = testData6[13045];
@(posedge clk);
#1;data_in = testData6[13046];
@(posedge clk);
#1;data_in = testData6[13047];
@(posedge clk);
#1;data_in = testData6[13048];
@(posedge clk);
#1;data_in = testData6[13049];
@(posedge clk);
#1;data_in = testData6[13050];
@(posedge clk);
#1;data_in = testData6[13051];
@(posedge clk);
#1;data_in = testData6[13052];
@(posedge clk);
#1;data_in = testData6[13053];
@(posedge clk);
#1;data_in = testData6[13054];
@(posedge clk);
#1;data_in = testData6[13055];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[13056];
@(posedge clk);
#1;data_in = testData6[13057];
@(posedge clk);
#1;data_in = testData6[13058];
@(posedge clk);
#1;data_in = testData6[13059];
@(posedge clk);
#1;data_in = testData6[13060];
@(posedge clk);
#1;data_in = testData6[13061];
@(posedge clk);
#1;data_in = testData6[13062];
@(posedge clk);
#1;data_in = testData6[13063];
@(posedge clk);
#1;data_in = testData6[13064];
@(posedge clk);
#1;data_in = testData6[13065];
@(posedge clk);
#1;data_in = testData6[13066];
@(posedge clk);
#1;data_in = testData6[13067];
@(posedge clk);
#1;data_in = testData6[13068];
@(posedge clk);
#1;data_in = testData6[13069];
@(posedge clk);
#1;data_in = testData6[13070];
@(posedge clk);
#1;data_in = testData6[13071];
@(posedge clk);
#1;data_in = testData6[13072];
@(posedge clk);
#1;data_in = testData6[13073];
@(posedge clk);
#1;data_in = testData6[13074];
@(posedge clk);
#1;data_in = testData6[13075];
@(posedge clk);
#1;data_in = testData6[13076];
@(posedge clk);
#1;data_in = testData6[13077];
@(posedge clk);
#1;data_in = testData6[13078];
@(posedge clk);
#1;data_in = testData6[13079];
@(posedge clk);
#1;data_in = testData6[13080];
@(posedge clk);
#1;data_in = testData6[13081];
@(posedge clk);
#1;data_in = testData6[13082];
@(posedge clk);
#1;data_in = testData6[13083];
@(posedge clk);
#1;data_in = testData6[13084];
@(posedge clk);
#1;data_in = testData6[13085];
@(posedge clk);
#1;data_in = testData6[13086];
@(posedge clk);
#1;data_in = testData6[13087];
@(posedge clk);
#1;data_in = testData6[13088];
@(posedge clk);
#1;data_in = testData6[13089];
@(posedge clk);
#1;data_in = testData6[13090];
@(posedge clk);
#1;data_in = testData6[13091];
@(posedge clk);
#1;data_in = testData6[13092];
@(posedge clk);
#1;data_in = testData6[13093];
@(posedge clk);
#1;data_in = testData6[13094];
@(posedge clk);
#1;data_in = testData6[13095];
@(posedge clk);
#1;data_in = testData6[13096];
@(posedge clk);
#1;data_in = testData6[13097];
@(posedge clk);
#1;data_in = testData6[13098];
@(posedge clk);
#1;data_in = testData6[13099];
@(posedge clk);
#1;data_in = testData6[13100];
@(posedge clk);
#1;data_in = testData6[13101];
@(posedge clk);
#1;data_in = testData6[13102];
@(posedge clk);
#1;data_in = testData6[13103];
@(posedge clk);
#1;data_in = testData6[13104];
@(posedge clk);
#1;data_in = testData6[13105];
@(posedge clk);
#1;data_in = testData6[13106];
@(posedge clk);
#1;data_in = testData6[13107];
@(posedge clk);
#1;data_in = testData6[13108];
@(posedge clk);
#1;data_in = testData6[13109];
@(posedge clk);
#1;data_in = testData6[13110];
@(posedge clk);
#1;data_in = testData6[13111];
@(posedge clk);
#1;data_in = testData6[13112];
@(posedge clk);
#1;data_in = testData6[13113];
@(posedge clk);
#1;data_in = testData6[13114];
@(posedge clk);
#1;data_in = testData6[13115];
@(posedge clk);
#1;data_in = testData6[13116];
@(posedge clk);
#1;data_in = testData6[13117];
@(posedge clk);
#1;data_in = testData6[13118];
@(posedge clk);
#1;data_in = testData6[13119];
@(posedge clk);
#1;data_in = testData6[13120];
@(posedge clk);
#1;data_in = testData6[13121];
@(posedge clk);
#1;data_in = testData6[13122];
@(posedge clk);
#1;data_in = testData6[13123];
@(posedge clk);
#1;data_in = testData6[13124];
@(posedge clk);
#1;data_in = testData6[13125];
@(posedge clk);
#1;data_in = testData6[13126];
@(posedge clk);
#1;data_in = testData6[13127];
@(posedge clk);
#1;data_in = testData6[13128];
@(posedge clk);
#1;data_in = testData6[13129];
@(posedge clk);
#1;data_in = testData6[13130];
@(posedge clk);
#1;data_in = testData6[13131];
@(posedge clk);
#1;data_in = testData6[13132];
@(posedge clk);
#1;data_in = testData6[13133];
@(posedge clk);
#1;data_in = testData6[13134];
@(posedge clk);
#1;data_in = testData6[13135];
@(posedge clk);
#1;data_in = testData6[13136];
@(posedge clk);
#1;data_in = testData6[13137];
@(posedge clk);
#1;data_in = testData6[13138];
@(posedge clk);
#1;data_in = testData6[13139];
@(posedge clk);
#1;data_in = testData6[13140];
@(posedge clk);
#1;data_in = testData6[13141];
@(posedge clk);
#1;data_in = testData6[13142];
@(posedge clk);
#1;data_in = testData6[13143];
@(posedge clk);
#1;data_in = testData6[13144];
@(posedge clk);
#1;data_in = testData6[13145];
@(posedge clk);
#1;data_in = testData6[13146];
@(posedge clk);
#1;data_in = testData6[13147];
@(posedge clk);
#1;data_in = testData6[13148];
@(posedge clk);
#1;data_in = testData6[13149];
@(posedge clk);
#1;data_in = testData6[13150];
@(posedge clk);
#1;data_in = testData6[13151];
@(posedge clk);
#1;data_in = testData6[13152];
@(posedge clk);
#1;data_in = testData6[13153];
@(posedge clk);
#1;data_in = testData6[13154];
@(posedge clk);
#1;data_in = testData6[13155];
@(posedge clk);
#1;data_in = testData6[13156];
@(posedge clk);
#1;data_in = testData6[13157];
@(posedge clk);
#1;data_in = testData6[13158];
@(posedge clk);
#1;data_in = testData6[13159];
@(posedge clk);
#1;data_in = testData6[13160];
@(posedge clk);
#1;data_in = testData6[13161];
@(posedge clk);
#1;data_in = testData6[13162];
@(posedge clk);
#1;data_in = testData6[13163];
@(posedge clk);
#1;data_in = testData6[13164];
@(posedge clk);
#1;data_in = testData6[13165];
@(posedge clk);
#1;data_in = testData6[13166];
@(posedge clk);
#1;data_in = testData6[13167];
@(posedge clk);
#1;data_in = testData6[13168];
@(posedge clk);
#1;data_in = testData6[13169];
@(posedge clk);
#1;data_in = testData6[13170];
@(posedge clk);
#1;data_in = testData6[13171];
@(posedge clk);
#1;data_in = testData6[13172];
@(posedge clk);
#1;data_in = testData6[13173];
@(posedge clk);
#1;data_in = testData6[13174];
@(posedge clk);
#1;data_in = testData6[13175];
@(posedge clk);
#1;data_in = testData6[13176];
@(posedge clk);
#1;data_in = testData6[13177];
@(posedge clk);
#1;data_in = testData6[13178];
@(posedge clk);
#1;data_in = testData6[13179];
@(posedge clk);
#1;data_in = testData6[13180];
@(posedge clk);
#1;data_in = testData6[13181];
@(posedge clk);
#1;data_in = testData6[13182];
@(posedge clk);
#1;data_in = testData6[13183];
@(posedge clk);
#1;data_in = testData6[13184];
@(posedge clk);
#1;data_in = testData6[13185];
@(posedge clk);
#1;data_in = testData6[13186];
@(posedge clk);
#1;data_in = testData6[13187];
@(posedge clk);
#1;data_in = testData6[13188];
@(posedge clk);
#1;data_in = testData6[13189];
@(posedge clk);
#1;data_in = testData6[13190];
@(posedge clk);
#1;data_in = testData6[13191];
@(posedge clk);
#1;data_in = testData6[13192];
@(posedge clk);
#1;data_in = testData6[13193];
@(posedge clk);
#1;data_in = testData6[13194];
@(posedge clk);
#1;data_in = testData6[13195];
@(posedge clk);
#1;data_in = testData6[13196];
@(posedge clk);
#1;data_in = testData6[13197];
@(posedge clk);
#1;data_in = testData6[13198];
@(posedge clk);
#1;data_in = testData6[13199];
@(posedge clk);
#1;data_in = testData6[13200];
@(posedge clk);
#1;data_in = testData6[13201];
@(posedge clk);
#1;data_in = testData6[13202];
@(posedge clk);
#1;data_in = testData6[13203];
@(posedge clk);
#1;data_in = testData6[13204];
@(posedge clk);
#1;data_in = testData6[13205];
@(posedge clk);
#1;data_in = testData6[13206];
@(posedge clk);
#1;data_in = testData6[13207];
@(posedge clk);
#1;data_in = testData6[13208];
@(posedge clk);
#1;data_in = testData6[13209];
@(posedge clk);
#1;data_in = testData6[13210];
@(posedge clk);
#1;data_in = testData6[13211];
@(posedge clk);
#1;data_in = testData6[13212];
@(posedge clk);
#1;data_in = testData6[13213];
@(posedge clk);
#1;data_in = testData6[13214];
@(posedge clk);
#1;data_in = testData6[13215];
@(posedge clk);
#1;data_in = testData6[13216];
@(posedge clk);
#1;data_in = testData6[13217];
@(posedge clk);
#1;data_in = testData6[13218];
@(posedge clk);
#1;data_in = testData6[13219];
@(posedge clk);
#1;data_in = testData6[13220];
@(posedge clk);
#1;data_in = testData6[13221];
@(posedge clk);
#1;data_in = testData6[13222];
@(posedge clk);
#1;data_in = testData6[13223];
@(posedge clk);
#1;data_in = testData6[13224];
@(posedge clk);
#1;data_in = testData6[13225];
@(posedge clk);
#1;data_in = testData6[13226];
@(posedge clk);
#1;data_in = testData6[13227];
@(posedge clk);
#1;data_in = testData6[13228];
@(posedge clk);
#1;data_in = testData6[13229];
@(posedge clk);
#1;data_in = testData6[13230];
@(posedge clk);
#1;data_in = testData6[13231];
@(posedge clk);
#1;data_in = testData6[13232];
@(posedge clk);
#1;data_in = testData6[13233];
@(posedge clk);
#1;data_in = testData6[13234];
@(posedge clk);
#1;data_in = testData6[13235];
@(posedge clk);
#1;data_in = testData6[13236];
@(posedge clk);
#1;data_in = testData6[13237];
@(posedge clk);
#1;data_in = testData6[13238];
@(posedge clk);
#1;data_in = testData6[13239];
@(posedge clk);
#1;data_in = testData6[13240];
@(posedge clk);
#1;data_in = testData6[13241];
@(posedge clk);
#1;data_in = testData6[13242];
@(posedge clk);
#1;data_in = testData6[13243];
@(posedge clk);
#1;data_in = testData6[13244];
@(posedge clk);
#1;data_in = testData6[13245];
@(posedge clk);
#1;data_in = testData6[13246];
@(posedge clk);
#1;data_in = testData6[13247];
@(posedge clk);
#1;data_in = testData6[13248];
@(posedge clk);
#1;data_in = testData6[13249];
@(posedge clk);
#1;data_in = testData6[13250];
@(posedge clk);
#1;data_in = testData6[13251];
@(posedge clk);
#1;data_in = testData6[13252];
@(posedge clk);
#1;data_in = testData6[13253];
@(posedge clk);
#1;data_in = testData6[13254];
@(posedge clk);
#1;data_in = testData6[13255];
@(posedge clk);
#1;data_in = testData6[13256];
@(posedge clk);
#1;data_in = testData6[13257];
@(posedge clk);
#1;data_in = testData6[13258];
@(posedge clk);
#1;data_in = testData6[13259];
@(posedge clk);
#1;data_in = testData6[13260];
@(posedge clk);
#1;data_in = testData6[13261];
@(posedge clk);
#1;data_in = testData6[13262];
@(posedge clk);
#1;data_in = testData6[13263];
@(posedge clk);
#1;data_in = testData6[13264];
@(posedge clk);
#1;data_in = testData6[13265];
@(posedge clk);
#1;data_in = testData6[13266];
@(posedge clk);
#1;data_in = testData6[13267];
@(posedge clk);
#1;data_in = testData6[13268];
@(posedge clk);
#1;data_in = testData6[13269];
@(posedge clk);
#1;data_in = testData6[13270];
@(posedge clk);
#1;data_in = testData6[13271];
@(posedge clk);
#1;data_in = testData6[13272];
@(posedge clk);
#1;data_in = testData6[13273];
@(posedge clk);
#1;data_in = testData6[13274];
@(posedge clk);
#1;data_in = testData6[13275];
@(posedge clk);
#1;data_in = testData6[13276];
@(posedge clk);
#1;data_in = testData6[13277];
@(posedge clk);
#1;data_in = testData6[13278];
@(posedge clk);
#1;data_in = testData6[13279];
@(posedge clk);
#1;data_in = testData6[13280];
@(posedge clk);
#1;data_in = testData6[13281];
@(posedge clk);
#1;data_in = testData6[13282];
@(posedge clk);
#1;data_in = testData6[13283];
@(posedge clk);
#1;data_in = testData6[13284];
@(posedge clk);
#1;data_in = testData6[13285];
@(posedge clk);
#1;data_in = testData6[13286];
@(posedge clk);
#1;data_in = testData6[13287];
@(posedge clk);
#1;data_in = testData6[13288];
@(posedge clk);
#1;data_in = testData6[13289];
@(posedge clk);
#1;data_in = testData6[13290];
@(posedge clk);
#1;data_in = testData6[13291];
@(posedge clk);
#1;data_in = testData6[13292];
@(posedge clk);
#1;data_in = testData6[13293];
@(posedge clk);
#1;data_in = testData6[13294];
@(posedge clk);
#1;data_in = testData6[13295];
@(posedge clk);
#1;data_in = testData6[13296];
@(posedge clk);
#1;data_in = testData6[13297];
@(posedge clk);
#1;data_in = testData6[13298];
@(posedge clk);
#1;data_in = testData6[13299];
@(posedge clk);
#1;data_in = testData6[13300];
@(posedge clk);
#1;data_in = testData6[13301];
@(posedge clk);
#1;data_in = testData6[13302];
@(posedge clk);
#1;data_in = testData6[13303];
@(posedge clk);
#1;data_in = testData6[13304];
@(posedge clk);
#1;data_in = testData6[13305];
@(posedge clk);
#1;data_in = testData6[13306];
@(posedge clk);
#1;data_in = testData6[13307];
@(posedge clk);
#1;data_in = testData6[13308];
@(posedge clk);
#1;data_in = testData6[13309];
@(posedge clk);
#1;data_in = testData6[13310];
@(posedge clk);
#1;data_in = testData6[13311];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[13312]; 
@(posedge clk);
#1;data_in = testData6[13313];
@(posedge clk);
#1;data_in = testData6[13314];
@(posedge clk);
#1;data_in = testData6[13315];
@(posedge clk);
#1;data_in = testData6[13316];
@(posedge clk);
#1;data_in = testData6[13317];
@(posedge clk);
#1;data_in = testData6[13318];
@(posedge clk);
#1;data_in = testData6[13319];
@(posedge clk);
#1;data_in = testData6[13320];
@(posedge clk);
#1;data_in = testData6[13321];
@(posedge clk);
#1;data_in = testData6[13322];
@(posedge clk);
#1;data_in = testData6[13323];
@(posedge clk);
#1;data_in = testData6[13324];
@(posedge clk);
#1;data_in = testData6[13325];
@(posedge clk);
#1;data_in = testData6[13326];
@(posedge clk);
#1;data_in = testData6[13327];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[13328];
@(posedge clk);
#1;data_in = testData6[13329];
@(posedge clk);
#1;data_in = testData6[13330];
@(posedge clk);
#1;data_in = testData6[13331];
@(posedge clk);
#1;data_in = testData6[13332];
@(posedge clk);
#1;data_in = testData6[13333];
@(posedge clk);
#1;data_in = testData6[13334];
@(posedge clk);
#1;data_in = testData6[13335];
@(posedge clk);
#1;data_in = testData6[13336];
@(posedge clk);
#1;data_in = testData6[13337];
@(posedge clk);
#1;data_in = testData6[13338];
@(posedge clk);
#1;data_in = testData6[13339];
@(posedge clk);
#1;data_in = testData6[13340];
@(posedge clk);
#1;data_in = testData6[13341];
@(posedge clk);
#1;data_in = testData6[13342];
@(posedge clk);
#1;data_in = testData6[13343];
@(posedge clk);
#1;data_in = testData6[13344];
@(posedge clk);
#1;data_in = testData6[13345];
@(posedge clk);
#1;data_in = testData6[13346];
@(posedge clk);
#1;data_in = testData6[13347];
@(posedge clk);
#1;data_in = testData6[13348];
@(posedge clk);
#1;data_in = testData6[13349];
@(posedge clk);
#1;data_in = testData6[13350];
@(posedge clk);
#1;data_in = testData6[13351];
@(posedge clk);
#1;data_in = testData6[13352];
@(posedge clk);
#1;data_in = testData6[13353];
@(posedge clk);
#1;data_in = testData6[13354];
@(posedge clk);
#1;data_in = testData6[13355];
@(posedge clk);
#1;data_in = testData6[13356];
@(posedge clk);
#1;data_in = testData6[13357];
@(posedge clk);
#1;data_in = testData6[13358];
@(posedge clk);
#1;data_in = testData6[13359];
@(posedge clk);
#1;data_in = testData6[13360];
@(posedge clk);
#1;data_in = testData6[13361];
@(posedge clk);
#1;data_in = testData6[13362];
@(posedge clk);
#1;data_in = testData6[13363];
@(posedge clk);
#1;data_in = testData6[13364];
@(posedge clk);
#1;data_in = testData6[13365];
@(posedge clk);
#1;data_in = testData6[13366];
@(posedge clk);
#1;data_in = testData6[13367];
@(posedge clk);
#1;data_in = testData6[13368];
@(posedge clk);
#1;data_in = testData6[13369];
@(posedge clk);
#1;data_in = testData6[13370];
@(posedge clk);
#1;data_in = testData6[13371];
@(posedge clk);
#1;data_in = testData6[13372];
@(posedge clk);
#1;data_in = testData6[13373];
@(posedge clk);
#1;data_in = testData6[13374];
@(posedge clk);
#1;data_in = testData6[13375];
@(posedge clk);
#1;data_in = testData6[13376];
@(posedge clk);
#1;data_in = testData6[13377];
@(posedge clk);
#1;data_in = testData6[13378];
@(posedge clk);
#1;data_in = testData6[13379];
@(posedge clk);
#1;data_in = testData6[13380];
@(posedge clk);
#1;data_in = testData6[13381];
@(posedge clk);
#1;data_in = testData6[13382];
@(posedge clk);
#1;data_in = testData6[13383];
@(posedge clk);
#1;data_in = testData6[13384];
@(posedge clk);
#1;data_in = testData6[13385];
@(posedge clk);
#1;data_in = testData6[13386];
@(posedge clk);
#1;data_in = testData6[13387];
@(posedge clk);
#1;data_in = testData6[13388];
@(posedge clk);
#1;data_in = testData6[13389];
@(posedge clk);
#1;data_in = testData6[13390];
@(posedge clk);
#1;data_in = testData6[13391];
@(posedge clk);
#1;data_in = testData6[13392];
@(posedge clk);
#1;data_in = testData6[13393];
@(posedge clk);
#1;data_in = testData6[13394];
@(posedge clk);
#1;data_in = testData6[13395];
@(posedge clk);
#1;data_in = testData6[13396];
@(posedge clk);
#1;data_in = testData6[13397];
@(posedge clk);
#1;data_in = testData6[13398];
@(posedge clk);
#1;data_in = testData6[13399];
@(posedge clk);
#1;data_in = testData6[13400];
@(posedge clk);
#1;data_in = testData6[13401];
@(posedge clk);
#1;data_in = testData6[13402];
@(posedge clk);
#1;data_in = testData6[13403];
@(posedge clk);
#1;data_in = testData6[13404];
@(posedge clk);
#1;data_in = testData6[13405];
@(posedge clk);
#1;data_in = testData6[13406];
@(posedge clk);
#1;data_in = testData6[13407];
@(posedge clk);
#1;data_in = testData6[13408];
@(posedge clk);
#1;data_in = testData6[13409];
@(posedge clk);
#1;data_in = testData6[13410];
@(posedge clk);
#1;data_in = testData6[13411];
@(posedge clk);
#1;data_in = testData6[13412];
@(posedge clk);
#1;data_in = testData6[13413];
@(posedge clk);
#1;data_in = testData6[13414];
@(posedge clk);
#1;data_in = testData6[13415];
@(posedge clk);
#1;data_in = testData6[13416];
@(posedge clk);
#1;data_in = testData6[13417];
@(posedge clk);
#1;data_in = testData6[13418];
@(posedge clk);
#1;data_in = testData6[13419];
@(posedge clk);
#1;data_in = testData6[13420];
@(posedge clk);
#1;data_in = testData6[13421];
@(posedge clk);
#1;data_in = testData6[13422];
@(posedge clk);
#1;data_in = testData6[13423];
@(posedge clk);
#1;data_in = testData6[13424];
@(posedge clk);
#1;data_in = testData6[13425];
@(posedge clk);
#1;data_in = testData6[13426];
@(posedge clk);
#1;data_in = testData6[13427];
@(posedge clk);
#1;data_in = testData6[13428];
@(posedge clk);
#1;data_in = testData6[13429];
@(posedge clk);
#1;data_in = testData6[13430];
@(posedge clk);
#1;data_in = testData6[13431];
@(posedge clk);
#1;data_in = testData6[13432];
@(posedge clk);
#1;data_in = testData6[13433];
@(posedge clk);
#1;data_in = testData6[13434];
@(posedge clk);
#1;data_in = testData6[13435];
@(posedge clk);
#1;data_in = testData6[13436];
@(posedge clk);
#1;data_in = testData6[13437];
@(posedge clk);
#1;data_in = testData6[13438];
@(posedge clk);
#1;data_in = testData6[13439];
@(posedge clk);
#1;data_in = testData6[13440];
@(posedge clk);
#1;data_in = testData6[13441];
@(posedge clk);
#1;data_in = testData6[13442];
@(posedge clk);
#1;data_in = testData6[13443];
@(posedge clk);
#1;data_in = testData6[13444];
@(posedge clk);
#1;data_in = testData6[13445];
@(posedge clk);
#1;data_in = testData6[13446];
@(posedge clk);
#1;data_in = testData6[13447];
@(posedge clk);
#1;data_in = testData6[13448];
@(posedge clk);
#1;data_in = testData6[13449];
@(posedge clk);
#1;data_in = testData6[13450];
@(posedge clk);
#1;data_in = testData6[13451];
@(posedge clk);
#1;data_in = testData6[13452];
@(posedge clk);
#1;data_in = testData6[13453];
@(posedge clk);
#1;data_in = testData6[13454];
@(posedge clk);
#1;data_in = testData6[13455];
@(posedge clk);
#1;data_in = testData6[13456];
@(posedge clk);
#1;data_in = testData6[13457];
@(posedge clk);
#1;data_in = testData6[13458];
@(posedge clk);
#1;data_in = testData6[13459];
@(posedge clk);
#1;data_in = testData6[13460];
@(posedge clk);
#1;data_in = testData6[13461];
@(posedge clk);
#1;data_in = testData6[13462];
@(posedge clk);
#1;data_in = testData6[13463];
@(posedge clk);
#1;data_in = testData6[13464];
@(posedge clk);
#1;data_in = testData6[13465];
@(posedge clk);
#1;data_in = testData6[13466];
@(posedge clk);
#1;data_in = testData6[13467];
@(posedge clk);
#1;data_in = testData6[13468];
@(posedge clk);
#1;data_in = testData6[13469];
@(posedge clk);
#1;data_in = testData6[13470];
@(posedge clk);
#1;data_in = testData6[13471];
@(posedge clk);
#1;data_in = testData6[13472];
@(posedge clk);
#1;data_in = testData6[13473];
@(posedge clk);
#1;data_in = testData6[13474];
@(posedge clk);
#1;data_in = testData6[13475];
@(posedge clk);
#1;data_in = testData6[13476];
@(posedge clk);
#1;data_in = testData6[13477];
@(posedge clk);
#1;data_in = testData6[13478];
@(posedge clk);
#1;data_in = testData6[13479];
@(posedge clk);
#1;data_in = testData6[13480];
@(posedge clk);
#1;data_in = testData6[13481];
@(posedge clk);
#1;data_in = testData6[13482];
@(posedge clk);
#1;data_in = testData6[13483];
@(posedge clk);
#1;data_in = testData6[13484];
@(posedge clk);
#1;data_in = testData6[13485];
@(posedge clk);
#1;data_in = testData6[13486];
@(posedge clk);
#1;data_in = testData6[13487];
@(posedge clk);
#1;data_in = testData6[13488];
@(posedge clk);
#1;data_in = testData6[13489];
@(posedge clk);
#1;data_in = testData6[13490];
@(posedge clk);
#1;data_in = testData6[13491];
@(posedge clk);
#1;data_in = testData6[13492];
@(posedge clk);
#1;data_in = testData6[13493];
@(posedge clk);
#1;data_in = testData6[13494];
@(posedge clk);
#1;data_in = testData6[13495];
@(posedge clk);
#1;data_in = testData6[13496];
@(posedge clk);
#1;data_in = testData6[13497];
@(posedge clk);
#1;data_in = testData6[13498];
@(posedge clk);
#1;data_in = testData6[13499];
@(posedge clk);
#1;data_in = testData6[13500];
@(posedge clk);
#1;data_in = testData6[13501];
@(posedge clk);
#1;data_in = testData6[13502];
@(posedge clk);
#1;data_in = testData6[13503];
@(posedge clk);
#1;data_in = testData6[13504];
@(posedge clk);
#1;data_in = testData6[13505];
@(posedge clk);
#1;data_in = testData6[13506];
@(posedge clk);
#1;data_in = testData6[13507];
@(posedge clk);
#1;data_in = testData6[13508];
@(posedge clk);
#1;data_in = testData6[13509];
@(posedge clk);
#1;data_in = testData6[13510];
@(posedge clk);
#1;data_in = testData6[13511];
@(posedge clk);
#1;data_in = testData6[13512];
@(posedge clk);
#1;data_in = testData6[13513];
@(posedge clk);
#1;data_in = testData6[13514];
@(posedge clk);
#1;data_in = testData6[13515];
@(posedge clk);
#1;data_in = testData6[13516];
@(posedge clk);
#1;data_in = testData6[13517];
@(posedge clk);
#1;data_in = testData6[13518];
@(posedge clk);
#1;data_in = testData6[13519];
@(posedge clk);
#1;data_in = testData6[13520];
@(posedge clk);
#1;data_in = testData6[13521];
@(posedge clk);
#1;data_in = testData6[13522];
@(posedge clk);
#1;data_in = testData6[13523];
@(posedge clk);
#1;data_in = testData6[13524];
@(posedge clk);
#1;data_in = testData6[13525];
@(posedge clk);
#1;data_in = testData6[13526];
@(posedge clk);
#1;data_in = testData6[13527];
@(posedge clk);
#1;data_in = testData6[13528];
@(posedge clk);
#1;data_in = testData6[13529];
@(posedge clk);
#1;data_in = testData6[13530];
@(posedge clk);
#1;data_in = testData6[13531];
@(posedge clk);
#1;data_in = testData6[13532];
@(posedge clk);
#1;data_in = testData6[13533];
@(posedge clk);
#1;data_in = testData6[13534];
@(posedge clk);
#1;data_in = testData6[13535];
@(posedge clk);
#1;data_in = testData6[13536];
@(posedge clk);
#1;data_in = testData6[13537];
@(posedge clk);
#1;data_in = testData6[13538];
@(posedge clk);
#1;data_in = testData6[13539];
@(posedge clk);
#1;data_in = testData6[13540];
@(posedge clk);
#1;data_in = testData6[13541];
@(posedge clk);
#1;data_in = testData6[13542];
@(posedge clk);
#1;data_in = testData6[13543];
@(posedge clk);
#1;data_in = testData6[13544];
@(posedge clk);
#1;data_in = testData6[13545];
@(posedge clk);
#1;data_in = testData6[13546];
@(posedge clk);
#1;data_in = testData6[13547];
@(posedge clk);
#1;data_in = testData6[13548];
@(posedge clk);
#1;data_in = testData6[13549];
@(posedge clk);
#1;data_in = testData6[13550];
@(posedge clk);
#1;data_in = testData6[13551];
@(posedge clk);
#1;data_in = testData6[13552];
@(posedge clk);
#1;data_in = testData6[13553];
@(posedge clk);
#1;data_in = testData6[13554];
@(posedge clk);
#1;data_in = testData6[13555];
@(posedge clk);
#1;data_in = testData6[13556];
@(posedge clk);
#1;data_in = testData6[13557];
@(posedge clk);
#1;data_in = testData6[13558];
@(posedge clk);
#1;data_in = testData6[13559];
@(posedge clk);
#1;data_in = testData6[13560];
@(posedge clk);
#1;data_in = testData6[13561];
@(posedge clk);
#1;data_in = testData6[13562];
@(posedge clk);
#1;data_in = testData6[13563];
@(posedge clk);
#1;data_in = testData6[13564];
@(posedge clk);
#1;data_in = testData6[13565];
@(posedge clk);
#1;data_in = testData6[13566];
@(posedge clk);
#1;data_in = testData6[13567];
@(posedge clk);
#1;data_in = testData6[13568];
@(posedge clk);
#1;data_in = testData6[13569];
@(posedge clk);
#1;data_in = testData6[13570];
@(posedge clk);
#1;data_in = testData6[13571];
@(posedge clk);
#1;data_in = testData6[13572];
@(posedge clk);
#1;data_in = testData6[13573];
@(posedge clk);
#1;data_in = testData6[13574];
@(posedge clk);
#1;data_in = testData6[13575];
@(posedge clk);
#1;data_in = testData6[13576];
@(posedge clk);
#1;data_in = testData6[13577];
@(posedge clk);
#1;data_in = testData6[13578];
@(posedge clk);
#1;data_in = testData6[13579];
@(posedge clk);
#1;data_in = testData6[13580];
@(posedge clk);
#1;data_in = testData6[13581];
@(posedge clk);
#1;data_in = testData6[13582];
@(posedge clk);
#1;data_in = testData6[13583];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[13584]; 
@(posedge clk);
#1;data_in = testData6[13585];
@(posedge clk);
#1;data_in = testData6[13586];
@(posedge clk);
#1;data_in = testData6[13587];
@(posedge clk);
#1;data_in = testData6[13588];
@(posedge clk);
#1;data_in = testData6[13589];
@(posedge clk);
#1;data_in = testData6[13590];
@(posedge clk);
#1;data_in = testData6[13591];
@(posedge clk);
#1;data_in = testData6[13592];
@(posedge clk);
#1;data_in = testData6[13593];
@(posedge clk);
#1;data_in = testData6[13594];
@(posedge clk);
#1;data_in = testData6[13595];
@(posedge clk);
#1;data_in = testData6[13596];
@(posedge clk);
#1;data_in = testData6[13597];
@(posedge clk);
#1;data_in = testData6[13598];
@(posedge clk);
#1;data_in = testData6[13599];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[13600];
@(posedge clk);
#1;data_in = testData6[13601];
@(posedge clk);
#1;data_in = testData6[13602];
@(posedge clk);
#1;data_in = testData6[13603];
@(posedge clk);
#1;data_in = testData6[13604];
@(posedge clk);
#1;data_in = testData6[13605];
@(posedge clk);
#1;data_in = testData6[13606];
@(posedge clk);
#1;data_in = testData6[13607];
@(posedge clk);
#1;data_in = testData6[13608];
@(posedge clk);
#1;data_in = testData6[13609];
@(posedge clk);
#1;data_in = testData6[13610];
@(posedge clk);
#1;data_in = testData6[13611];
@(posedge clk);
#1;data_in = testData6[13612];
@(posedge clk);
#1;data_in = testData6[13613];
@(posedge clk);
#1;data_in = testData6[13614];
@(posedge clk);
#1;data_in = testData6[13615];
@(posedge clk);
#1;data_in = testData6[13616];
@(posedge clk);
#1;data_in = testData6[13617];
@(posedge clk);
#1;data_in = testData6[13618];
@(posedge clk);
#1;data_in = testData6[13619];
@(posedge clk);
#1;data_in = testData6[13620];
@(posedge clk);
#1;data_in = testData6[13621];
@(posedge clk);
#1;data_in = testData6[13622];
@(posedge clk);
#1;data_in = testData6[13623];
@(posedge clk);
#1;data_in = testData6[13624];
@(posedge clk);
#1;data_in = testData6[13625];
@(posedge clk);
#1;data_in = testData6[13626];
@(posedge clk);
#1;data_in = testData6[13627];
@(posedge clk);
#1;data_in = testData6[13628];
@(posedge clk);
#1;data_in = testData6[13629];
@(posedge clk);
#1;data_in = testData6[13630];
@(posedge clk);
#1;data_in = testData6[13631];
@(posedge clk);
#1;data_in = testData6[13632];
@(posedge clk);
#1;data_in = testData6[13633];
@(posedge clk);
#1;data_in = testData6[13634];
@(posedge clk);
#1;data_in = testData6[13635];
@(posedge clk);
#1;data_in = testData6[13636];
@(posedge clk);
#1;data_in = testData6[13637];
@(posedge clk);
#1;data_in = testData6[13638];
@(posedge clk);
#1;data_in = testData6[13639];
@(posedge clk);
#1;data_in = testData6[13640];
@(posedge clk);
#1;data_in = testData6[13641];
@(posedge clk);
#1;data_in = testData6[13642];
@(posedge clk);
#1;data_in = testData6[13643];
@(posedge clk);
#1;data_in = testData6[13644];
@(posedge clk);
#1;data_in = testData6[13645];
@(posedge clk);
#1;data_in = testData6[13646];
@(posedge clk);
#1;data_in = testData6[13647];
@(posedge clk);
#1;data_in = testData6[13648];
@(posedge clk);
#1;data_in = testData6[13649];
@(posedge clk);
#1;data_in = testData6[13650];
@(posedge clk);
#1;data_in = testData6[13651];
@(posedge clk);
#1;data_in = testData6[13652];
@(posedge clk);
#1;data_in = testData6[13653];
@(posedge clk);
#1;data_in = testData6[13654];
@(posedge clk);
#1;data_in = testData6[13655];
@(posedge clk);
#1;data_in = testData6[13656];
@(posedge clk);
#1;data_in = testData6[13657];
@(posedge clk);
#1;data_in = testData6[13658];
@(posedge clk);
#1;data_in = testData6[13659];
@(posedge clk);
#1;data_in = testData6[13660];
@(posedge clk);
#1;data_in = testData6[13661];
@(posedge clk);
#1;data_in = testData6[13662];
@(posedge clk);
#1;data_in = testData6[13663];
@(posedge clk);
#1;data_in = testData6[13664];
@(posedge clk);
#1;data_in = testData6[13665];
@(posedge clk);
#1;data_in = testData6[13666];
@(posedge clk);
#1;data_in = testData6[13667];
@(posedge clk);
#1;data_in = testData6[13668];
@(posedge clk);
#1;data_in = testData6[13669];
@(posedge clk);
#1;data_in = testData6[13670];
@(posedge clk);
#1;data_in = testData6[13671];
@(posedge clk);
#1;data_in = testData6[13672];
@(posedge clk);
#1;data_in = testData6[13673];
@(posedge clk);
#1;data_in = testData6[13674];
@(posedge clk);
#1;data_in = testData6[13675];
@(posedge clk);
#1;data_in = testData6[13676];
@(posedge clk);
#1;data_in = testData6[13677];
@(posedge clk);
#1;data_in = testData6[13678];
@(posedge clk);
#1;data_in = testData6[13679];
@(posedge clk);
#1;data_in = testData6[13680];
@(posedge clk);
#1;data_in = testData6[13681];
@(posedge clk);
#1;data_in = testData6[13682];
@(posedge clk);
#1;data_in = testData6[13683];
@(posedge clk);
#1;data_in = testData6[13684];
@(posedge clk);
#1;data_in = testData6[13685];
@(posedge clk);
#1;data_in = testData6[13686];
@(posedge clk);
#1;data_in = testData6[13687];
@(posedge clk);
#1;data_in = testData6[13688];
@(posedge clk);
#1;data_in = testData6[13689];
@(posedge clk);
#1;data_in = testData6[13690];
@(posedge clk);
#1;data_in = testData6[13691];
@(posedge clk);
#1;data_in = testData6[13692];
@(posedge clk);
#1;data_in = testData6[13693];
@(posedge clk);
#1;data_in = testData6[13694];
@(posedge clk);
#1;data_in = testData6[13695];
@(posedge clk);
#1;data_in = testData6[13696];
@(posedge clk);
#1;data_in = testData6[13697];
@(posedge clk);
#1;data_in = testData6[13698];
@(posedge clk);
#1;data_in = testData6[13699];
@(posedge clk);
#1;data_in = testData6[13700];
@(posedge clk);
#1;data_in = testData6[13701];
@(posedge clk);
#1;data_in = testData6[13702];
@(posedge clk);
#1;data_in = testData6[13703];
@(posedge clk);
#1;data_in = testData6[13704];
@(posedge clk);
#1;data_in = testData6[13705];
@(posedge clk);
#1;data_in = testData6[13706];
@(posedge clk);
#1;data_in = testData6[13707];
@(posedge clk);
#1;data_in = testData6[13708];
@(posedge clk);
#1;data_in = testData6[13709];
@(posedge clk);
#1;data_in = testData6[13710];
@(posedge clk);
#1;data_in = testData6[13711];
@(posedge clk);
#1;data_in = testData6[13712];
@(posedge clk);
#1;data_in = testData6[13713];
@(posedge clk);
#1;data_in = testData6[13714];
@(posedge clk);
#1;data_in = testData6[13715];
@(posedge clk);
#1;data_in = testData6[13716];
@(posedge clk);
#1;data_in = testData6[13717];
@(posedge clk);
#1;data_in = testData6[13718];
@(posedge clk);
#1;data_in = testData6[13719];
@(posedge clk);
#1;data_in = testData6[13720];
@(posedge clk);
#1;data_in = testData6[13721];
@(posedge clk);
#1;data_in = testData6[13722];
@(posedge clk);
#1;data_in = testData6[13723];
@(posedge clk);
#1;data_in = testData6[13724];
@(posedge clk);
#1;data_in = testData6[13725];
@(posedge clk);
#1;data_in = testData6[13726];
@(posedge clk);
#1;data_in = testData6[13727];
@(posedge clk);
#1;data_in = testData6[13728];
@(posedge clk);
#1;data_in = testData6[13729];
@(posedge clk);
#1;data_in = testData6[13730];
@(posedge clk);
#1;data_in = testData6[13731];
@(posedge clk);
#1;data_in = testData6[13732];
@(posedge clk);
#1;data_in = testData6[13733];
@(posedge clk);
#1;data_in = testData6[13734];
@(posedge clk);
#1;data_in = testData6[13735];
@(posedge clk);
#1;data_in = testData6[13736];
@(posedge clk);
#1;data_in = testData6[13737];
@(posedge clk);
#1;data_in = testData6[13738];
@(posedge clk);
#1;data_in = testData6[13739];
@(posedge clk);
#1;data_in = testData6[13740];
@(posedge clk);
#1;data_in = testData6[13741];
@(posedge clk);
#1;data_in = testData6[13742];
@(posedge clk);
#1;data_in = testData6[13743];
@(posedge clk);
#1;data_in = testData6[13744];
@(posedge clk);
#1;data_in = testData6[13745];
@(posedge clk);
#1;data_in = testData6[13746];
@(posedge clk);
#1;data_in = testData6[13747];
@(posedge clk);
#1;data_in = testData6[13748];
@(posedge clk);
#1;data_in = testData6[13749];
@(posedge clk);
#1;data_in = testData6[13750];
@(posedge clk);
#1;data_in = testData6[13751];
@(posedge clk);
#1;data_in = testData6[13752];
@(posedge clk);
#1;data_in = testData6[13753];
@(posedge clk);
#1;data_in = testData6[13754];
@(posedge clk);
#1;data_in = testData6[13755];
@(posedge clk);
#1;data_in = testData6[13756];
@(posedge clk);
#1;data_in = testData6[13757];
@(posedge clk);
#1;data_in = testData6[13758];
@(posedge clk);
#1;data_in = testData6[13759];
@(posedge clk);
#1;data_in = testData6[13760];
@(posedge clk);
#1;data_in = testData6[13761];
@(posedge clk);
#1;data_in = testData6[13762];
@(posedge clk);
#1;data_in = testData6[13763];
@(posedge clk);
#1;data_in = testData6[13764];
@(posedge clk);
#1;data_in = testData6[13765];
@(posedge clk);
#1;data_in = testData6[13766];
@(posedge clk);
#1;data_in = testData6[13767];
@(posedge clk);
#1;data_in = testData6[13768];
@(posedge clk);
#1;data_in = testData6[13769];
@(posedge clk);
#1;data_in = testData6[13770];
@(posedge clk);
#1;data_in = testData6[13771];
@(posedge clk);
#1;data_in = testData6[13772];
@(posedge clk);
#1;data_in = testData6[13773];
@(posedge clk);
#1;data_in = testData6[13774];
@(posedge clk);
#1;data_in = testData6[13775];
@(posedge clk);
#1;data_in = testData6[13776];
@(posedge clk);
#1;data_in = testData6[13777];
@(posedge clk);
#1;data_in = testData6[13778];
@(posedge clk);
#1;data_in = testData6[13779];
@(posedge clk);
#1;data_in = testData6[13780];
@(posedge clk);
#1;data_in = testData6[13781];
@(posedge clk);
#1;data_in = testData6[13782];
@(posedge clk);
#1;data_in = testData6[13783];
@(posedge clk);
#1;data_in = testData6[13784];
@(posedge clk);
#1;data_in = testData6[13785];
@(posedge clk);
#1;data_in = testData6[13786];
@(posedge clk);
#1;data_in = testData6[13787];
@(posedge clk);
#1;data_in = testData6[13788];
@(posedge clk);
#1;data_in = testData6[13789];
@(posedge clk);
#1;data_in = testData6[13790];
@(posedge clk);
#1;data_in = testData6[13791];
@(posedge clk);
#1;data_in = testData6[13792];
@(posedge clk);
#1;data_in = testData6[13793];
@(posedge clk);
#1;data_in = testData6[13794];
@(posedge clk);
#1;data_in = testData6[13795];
@(posedge clk);
#1;data_in = testData6[13796];
@(posedge clk);
#1;data_in = testData6[13797];
@(posedge clk);
#1;data_in = testData6[13798];
@(posedge clk);
#1;data_in = testData6[13799];
@(posedge clk);
#1;data_in = testData6[13800];
@(posedge clk);
#1;data_in = testData6[13801];
@(posedge clk);
#1;data_in = testData6[13802];
@(posedge clk);
#1;data_in = testData6[13803];
@(posedge clk);
#1;data_in = testData6[13804];
@(posedge clk);
#1;data_in = testData6[13805];
@(posedge clk);
#1;data_in = testData6[13806];
@(posedge clk);
#1;data_in = testData6[13807];
@(posedge clk);
#1;data_in = testData6[13808];
@(posedge clk);
#1;data_in = testData6[13809];
@(posedge clk);
#1;data_in = testData6[13810];
@(posedge clk);
#1;data_in = testData6[13811];
@(posedge clk);
#1;data_in = testData6[13812];
@(posedge clk);
#1;data_in = testData6[13813];
@(posedge clk);
#1;data_in = testData6[13814];
@(posedge clk);
#1;data_in = testData6[13815];
@(posedge clk);
#1;data_in = testData6[13816];
@(posedge clk);
#1;data_in = testData6[13817];
@(posedge clk);
#1;data_in = testData6[13818];
@(posedge clk);
#1;data_in = testData6[13819];
@(posedge clk);
#1;data_in = testData6[13820];
@(posedge clk);
#1;data_in = testData6[13821];
@(posedge clk);
#1;data_in = testData6[13822];
@(posedge clk);
#1;data_in = testData6[13823];
@(posedge clk);
#1;data_in = testData6[13824];
@(posedge clk);
#1;data_in = testData6[13825];
@(posedge clk);
#1;data_in = testData6[13826];
@(posedge clk);
#1;data_in = testData6[13827];
@(posedge clk);
#1;data_in = testData6[13828];
@(posedge clk);
#1;data_in = testData6[13829];
@(posedge clk);
#1;data_in = testData6[13830];
@(posedge clk);
#1;data_in = testData6[13831];
@(posedge clk);
#1;data_in = testData6[13832];
@(posedge clk);
#1;data_in = testData6[13833];
@(posedge clk);
#1;data_in = testData6[13834];
@(posedge clk);
#1;data_in = testData6[13835];
@(posedge clk);
#1;data_in = testData6[13836];
@(posedge clk);
#1;data_in = testData6[13837];
@(posedge clk);
#1;data_in = testData6[13838];
@(posedge clk);
#1;data_in = testData6[13839];
@(posedge clk);
#1;data_in = testData6[13840];
@(posedge clk);
#1;data_in = testData6[13841];
@(posedge clk);
#1;data_in = testData6[13842];
@(posedge clk);
#1;data_in = testData6[13843];
@(posedge clk);
#1;data_in = testData6[13844];
@(posedge clk);
#1;data_in = testData6[13845];
@(posedge clk);
#1;data_in = testData6[13846];
@(posedge clk);
#1;data_in = testData6[13847];
@(posedge clk);
#1;data_in = testData6[13848];
@(posedge clk);
#1;data_in = testData6[13849];
@(posedge clk);
#1;data_in = testData6[13850];
@(posedge clk);
#1;data_in = testData6[13851];
@(posedge clk);
#1;data_in = testData6[13852];
@(posedge clk);
#1;data_in = testData6[13853];
@(posedge clk);
#1;data_in = testData6[13854];
@(posedge clk);
#1;data_in = testData6[13855];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[13856]; 
@(posedge clk);
#1;data_in = testData6[13857];
@(posedge clk);
#1;data_in = testData6[13858];
@(posedge clk);
#1;data_in = testData6[13859];
@(posedge clk);
#1;data_in = testData6[13860];
@(posedge clk);
#1;data_in = testData6[13861];
@(posedge clk);
#1;data_in = testData6[13862];
@(posedge clk);
#1;data_in = testData6[13863];
@(posedge clk);
#1;data_in = testData6[13864];
@(posedge clk);
#1;data_in = testData6[13865];
@(posedge clk);
#1;data_in = testData6[13866];
@(posedge clk);
#1;data_in = testData6[13867];
@(posedge clk);
#1;data_in = testData6[13868];
@(posedge clk);
#1;data_in = testData6[13869];
@(posedge clk);
#1;data_in = testData6[13870];
@(posedge clk);
#1;data_in = testData6[13871];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=16, p=16, b=8, g=1

module tb5();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_16_16_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData5[13071:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb5", testData5);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb5");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData5[0];
@(posedge clk);
#1;data_in = testData5[1];
@(posedge clk);
#1;data_in = testData5[2];
@(posedge clk);
#1;data_in = testData5[3];
@(posedge clk);
#1;data_in = testData5[4];
@(posedge clk);
#1;data_in = testData5[5];
@(posedge clk);
#1;data_in = testData5[6];
@(posedge clk);
#1;data_in = testData5[7];
@(posedge clk);
#1;data_in = testData5[8];
@(posedge clk);
#1;data_in = testData5[9];
@(posedge clk);
#1;data_in = testData5[10];
@(posedge clk);
#1;data_in = testData5[11];
@(posedge clk);
#1;data_in = testData5[12];
@(posedge clk);
#1;data_in = testData5[13];
@(posedge clk);
#1;data_in = testData5[14];
@(posedge clk);
#1;data_in = testData5[15];
@(posedge clk);
#1;data_in = testData5[16];
@(posedge clk);
#1;data_in = testData5[17];
@(posedge clk);
#1;data_in = testData5[18];
@(posedge clk);
#1;data_in = testData5[19];
@(posedge clk);
#1;data_in = testData5[20];
@(posedge clk);
#1;data_in = testData5[21];
@(posedge clk);
#1;data_in = testData5[22];
@(posedge clk);
#1;data_in = testData5[23];
@(posedge clk);
#1;data_in = testData5[24];
@(posedge clk);
#1;data_in = testData5[25];
@(posedge clk);
#1;data_in = testData5[26];
@(posedge clk);
#1;data_in = testData5[27];
@(posedge clk);
#1;data_in = testData5[28];
@(posedge clk);
#1;data_in = testData5[29];
@(posedge clk);
#1;data_in = testData5[30];
@(posedge clk);
#1;data_in = testData5[31];
@(posedge clk);
#1;data_in = testData5[32];
@(posedge clk);
#1;data_in = testData5[33];
@(posedge clk);
#1;data_in = testData5[34];
@(posedge clk);
#1;data_in = testData5[35];
@(posedge clk);
#1;data_in = testData5[36];
@(posedge clk);
#1;data_in = testData5[37];
@(posedge clk);
#1;data_in = testData5[38];
@(posedge clk);
#1;data_in = testData5[39];
@(posedge clk);
#1;data_in = testData5[40];
@(posedge clk);
#1;data_in = testData5[41];
@(posedge clk);
#1;data_in = testData5[42];
@(posedge clk);
#1;data_in = testData5[43];
@(posedge clk);
#1;data_in = testData5[44];
@(posedge clk);
#1;data_in = testData5[45];
@(posedge clk);
#1;data_in = testData5[46];
@(posedge clk);
#1;data_in = testData5[47];
@(posedge clk);
#1;data_in = testData5[48];
@(posedge clk);
#1;data_in = testData5[49];
@(posedge clk);
#1;data_in = testData5[50];
@(posedge clk);
#1;data_in = testData5[51];
@(posedge clk);
#1;data_in = testData5[52];
@(posedge clk);
#1;data_in = testData5[53];
@(posedge clk);
#1;data_in = testData5[54];
@(posedge clk);
#1;data_in = testData5[55];
@(posedge clk);
#1;data_in = testData5[56];
@(posedge clk);
#1;data_in = testData5[57];
@(posedge clk);
#1;data_in = testData5[58];
@(posedge clk);
#1;data_in = testData5[59];
@(posedge clk);
#1;data_in = testData5[60];
@(posedge clk);
#1;data_in = testData5[61];
@(posedge clk);
#1;data_in = testData5[62];
@(posedge clk);
#1;data_in = testData5[63];
@(posedge clk);
#1;data_in = testData5[64];
@(posedge clk);
#1;data_in = testData5[65];
@(posedge clk);
#1;data_in = testData5[66];
@(posedge clk);
#1;data_in = testData5[67];
@(posedge clk);
#1;data_in = testData5[68];
@(posedge clk);
#1;data_in = testData5[69];
@(posedge clk);
#1;data_in = testData5[70];
@(posedge clk);
#1;data_in = testData5[71];
@(posedge clk);
#1;data_in = testData5[72];
@(posedge clk);
#1;data_in = testData5[73];
@(posedge clk);
#1;data_in = testData5[74];
@(posedge clk);
#1;data_in = testData5[75];
@(posedge clk);
#1;data_in = testData5[76];
@(posedge clk);
#1;data_in = testData5[77];
@(posedge clk);
#1;data_in = testData5[78];
@(posedge clk);
#1;data_in = testData5[79];
@(posedge clk);
#1;data_in = testData5[80];
@(posedge clk);
#1;data_in = testData5[81];
@(posedge clk);
#1;data_in = testData5[82];
@(posedge clk);
#1;data_in = testData5[83];
@(posedge clk);
#1;data_in = testData5[84];
@(posedge clk);
#1;data_in = testData5[85];
@(posedge clk);
#1;data_in = testData5[86];
@(posedge clk);
#1;data_in = testData5[87];
@(posedge clk);
#1;data_in = testData5[88];
@(posedge clk);
#1;data_in = testData5[89];
@(posedge clk);
#1;data_in = testData5[90];
@(posedge clk);
#1;data_in = testData5[91];
@(posedge clk);
#1;data_in = testData5[92];
@(posedge clk);
#1;data_in = testData5[93];
@(posedge clk);
#1;data_in = testData5[94];
@(posedge clk);
#1;data_in = testData5[95];
@(posedge clk);
#1;data_in = testData5[96];
@(posedge clk);
#1;data_in = testData5[97];
@(posedge clk);
#1;data_in = testData5[98];
@(posedge clk);
#1;data_in = testData5[99];
@(posedge clk);
#1;data_in = testData5[100];
@(posedge clk);
#1;data_in = testData5[101];
@(posedge clk);
#1;data_in = testData5[102];
@(posedge clk);
#1;data_in = testData5[103];
@(posedge clk);
#1;data_in = testData5[104];
@(posedge clk);
#1;data_in = testData5[105];
@(posedge clk);
#1;data_in = testData5[106];
@(posedge clk);
#1;data_in = testData5[107];
@(posedge clk);
#1;data_in = testData5[108];
@(posedge clk);
#1;data_in = testData5[109];
@(posedge clk);
#1;data_in = testData5[110];
@(posedge clk);
#1;data_in = testData5[111];
@(posedge clk);
#1;data_in = testData5[112];
@(posedge clk);
#1;data_in = testData5[113];
@(posedge clk);
#1;data_in = testData5[114];
@(posedge clk);
#1;data_in = testData5[115];
@(posedge clk);
#1;data_in = testData5[116];
@(posedge clk);
#1;data_in = testData5[117];
@(posedge clk);
#1;data_in = testData5[118];
@(posedge clk);
#1;data_in = testData5[119];
@(posedge clk);
#1;data_in = testData5[120];
@(posedge clk);
#1;data_in = testData5[121];
@(posedge clk);
#1;data_in = testData5[122];
@(posedge clk);
#1;data_in = testData5[123];
@(posedge clk);
#1;data_in = testData5[124];
@(posedge clk);
#1;data_in = testData5[125];
@(posedge clk);
#1;data_in = testData5[126];
@(posedge clk);
#1;data_in = testData5[127];
@(posedge clk);
#1;data_in = testData5[128];
@(posedge clk);
#1;data_in = testData5[129];
@(posedge clk);
#1;data_in = testData5[130];
@(posedge clk);
#1;data_in = testData5[131];
@(posedge clk);
#1;data_in = testData5[132];
@(posedge clk);
#1;data_in = testData5[133];
@(posedge clk);
#1;data_in = testData5[134];
@(posedge clk);
#1;data_in = testData5[135];
@(posedge clk);
#1;data_in = testData5[136];
@(posedge clk);
#1;data_in = testData5[137];
@(posedge clk);
#1;data_in = testData5[138];
@(posedge clk);
#1;data_in = testData5[139];
@(posedge clk);
#1;data_in = testData5[140];
@(posedge clk);
#1;data_in = testData5[141];
@(posedge clk);
#1;data_in = testData5[142];
@(posedge clk);
#1;data_in = testData5[143];
@(posedge clk);
#1;data_in = testData5[144];
@(posedge clk);
#1;data_in = testData5[145];
@(posedge clk);
#1;data_in = testData5[146];
@(posedge clk);
#1;data_in = testData5[147];
@(posedge clk);
#1;data_in = testData5[148];
@(posedge clk);
#1;data_in = testData5[149];
@(posedge clk);
#1;data_in = testData5[150];
@(posedge clk);
#1;data_in = testData5[151];
@(posedge clk);
#1;data_in = testData5[152];
@(posedge clk);
#1;data_in = testData5[153];
@(posedge clk);
#1;data_in = testData5[154];
@(posedge clk);
#1;data_in = testData5[155];
@(posedge clk);
#1;data_in = testData5[156];
@(posedge clk);
#1;data_in = testData5[157];
@(posedge clk);
#1;data_in = testData5[158];
@(posedge clk);
#1;data_in = testData5[159];
@(posedge clk);
#1;data_in = testData5[160];
@(posedge clk);
#1;data_in = testData5[161];
@(posedge clk);
#1;data_in = testData5[162];
@(posedge clk);
#1;data_in = testData5[163];
@(posedge clk);
#1;data_in = testData5[164];
@(posedge clk);
#1;data_in = testData5[165];
@(posedge clk);
#1;data_in = testData5[166];
@(posedge clk);
#1;data_in = testData5[167];
@(posedge clk);
#1;data_in = testData5[168];
@(posedge clk);
#1;data_in = testData5[169];
@(posedge clk);
#1;data_in = testData5[170];
@(posedge clk);
#1;data_in = testData5[171];
@(posedge clk);
#1;data_in = testData5[172];
@(posedge clk);
#1;data_in = testData5[173];
@(posedge clk);
#1;data_in = testData5[174];
@(posedge clk);
#1;data_in = testData5[175];
@(posedge clk);
#1;data_in = testData5[176];
@(posedge clk);
#1;data_in = testData5[177];
@(posedge clk);
#1;data_in = testData5[178];
@(posedge clk);
#1;data_in = testData5[179];
@(posedge clk);
#1;data_in = testData5[180];
@(posedge clk);
#1;data_in = testData5[181];
@(posedge clk);
#1;data_in = testData5[182];
@(posedge clk);
#1;data_in = testData5[183];
@(posedge clk);
#1;data_in = testData5[184];
@(posedge clk);
#1;data_in = testData5[185];
@(posedge clk);
#1;data_in = testData5[186];
@(posedge clk);
#1;data_in = testData5[187];
@(posedge clk);
#1;data_in = testData5[188];
@(posedge clk);
#1;data_in = testData5[189];
@(posedge clk);
#1;data_in = testData5[190];
@(posedge clk);
#1;data_in = testData5[191];
@(posedge clk);
#1;data_in = testData5[192];
@(posedge clk);
#1;data_in = testData5[193];
@(posedge clk);
#1;data_in = testData5[194];
@(posedge clk);
#1;data_in = testData5[195];
@(posedge clk);
#1;data_in = testData5[196];
@(posedge clk);
#1;data_in = testData5[197];
@(posedge clk);
#1;data_in = testData5[198];
@(posedge clk);
#1;data_in = testData5[199];
@(posedge clk);
#1;data_in = testData5[200];
@(posedge clk);
#1;data_in = testData5[201];
@(posedge clk);
#1;data_in = testData5[202];
@(posedge clk);
#1;data_in = testData5[203];
@(posedge clk);
#1;data_in = testData5[204];
@(posedge clk);
#1;data_in = testData5[205];
@(posedge clk);
#1;data_in = testData5[206];
@(posedge clk);
#1;data_in = testData5[207];
@(posedge clk);
#1;data_in = testData5[208];
@(posedge clk);
#1;data_in = testData5[209];
@(posedge clk);
#1;data_in = testData5[210];
@(posedge clk);
#1;data_in = testData5[211];
@(posedge clk);
#1;data_in = testData5[212];
@(posedge clk);
#1;data_in = testData5[213];
@(posedge clk);
#1;data_in = testData5[214];
@(posedge clk);
#1;data_in = testData5[215];
@(posedge clk);
#1;data_in = testData5[216];
@(posedge clk);
#1;data_in = testData5[217];
@(posedge clk);
#1;data_in = testData5[218];
@(posedge clk);
#1;data_in = testData5[219];
@(posedge clk);
#1;data_in = testData5[220];
@(posedge clk);
#1;data_in = testData5[221];
@(posedge clk);
#1;data_in = testData5[222];
@(posedge clk);
#1;data_in = testData5[223];
@(posedge clk);
#1;data_in = testData5[224];
@(posedge clk);
#1;data_in = testData5[225];
@(posedge clk);
#1;data_in = testData5[226];
@(posedge clk);
#1;data_in = testData5[227];
@(posedge clk);
#1;data_in = testData5[228];
@(posedge clk);
#1;data_in = testData5[229];
@(posedge clk);
#1;data_in = testData5[230];
@(posedge clk);
#1;data_in = testData5[231];
@(posedge clk);
#1;data_in = testData5[232];
@(posedge clk);
#1;data_in = testData5[233];
@(posedge clk);
#1;data_in = testData5[234];
@(posedge clk);
#1;data_in = testData5[235];
@(posedge clk);
#1;data_in = testData5[236];
@(posedge clk);
#1;data_in = testData5[237];
@(posedge clk);
#1;data_in = testData5[238];
@(posedge clk);
#1;data_in = testData5[239];
@(posedge clk);
#1;data_in = testData5[240];
@(posedge clk);
#1;data_in = testData5[241];
@(posedge clk);
#1;data_in = testData5[242];
@(posedge clk);
#1;data_in = testData5[243];
@(posedge clk);
#1;data_in = testData5[244];
@(posedge clk);
#1;data_in = testData5[245];
@(posedge clk);
#1;data_in = testData5[246];
@(posedge clk);
#1;data_in = testData5[247];
@(posedge clk);
#1;data_in = testData5[248];
@(posedge clk);
#1;data_in = testData5[249];
@(posedge clk);
#1;data_in = testData5[250];
@(posedge clk);
#1;data_in = testData5[251];
@(posedge clk);
#1;data_in = testData5[252];
@(posedge clk);
#1;data_in = testData5[253];
@(posedge clk);
#1;data_in = testData5[254];
@(posedge clk);
#1;data_in = testData5[255];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData5[256]; 
@(posedge clk);
#1;data_in = testData5[257];
@(posedge clk);
#1;data_in = testData5[258];
@(posedge clk);
#1;data_in = testData5[259];
@(posedge clk);
#1;data_in = testData5[260];
@(posedge clk);
#1;data_in = testData5[261];
@(posedge clk);
#1;data_in = testData5[262];
@(posedge clk);
#1;data_in = testData5[263];
@(posedge clk);
#1;data_in = testData5[264];
@(posedge clk);
#1;data_in = testData5[265];
@(posedge clk);
#1;data_in = testData5[266];
@(posedge clk);
#1;data_in = testData5[267];
@(posedge clk);
#1;data_in = testData5[268];
@(posedge clk);
#1;data_in = testData5[269];
@(posedge clk);
#1;data_in = testData5[270];
@(posedge clk);
#1;data_in = testData5[271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[272]; 
@(posedge clk);
#1;data_in = testData5[273];
@(posedge clk);
#1;data_in = testData5[274];
@(posedge clk);
#1;data_in = testData5[275];
@(posedge clk);
#1;data_in = testData5[276];
@(posedge clk);
#1;data_in = testData5[277];
@(posedge clk);
#1;data_in = testData5[278];
@(posedge clk);
#1;data_in = testData5[279];
@(posedge clk);
#1;data_in = testData5[280];
@(posedge clk);
#1;data_in = testData5[281];
@(posedge clk);
#1;data_in = testData5[282];
@(posedge clk);
#1;data_in = testData5[283];
@(posedge clk);
#1;data_in = testData5[284];
@(posedge clk);
#1;data_in = testData5[285];
@(posedge clk);
#1;data_in = testData5[286];
@(posedge clk);
#1;data_in = testData5[287];
@(posedge clk);
#1;data_in = testData5[288];
@(posedge clk);
#1;data_in = testData5[289];
@(posedge clk);
#1;data_in = testData5[290];
@(posedge clk);
#1;data_in = testData5[291];
@(posedge clk);
#1;data_in = testData5[292];
@(posedge clk);
#1;data_in = testData5[293];
@(posedge clk);
#1;data_in = testData5[294];
@(posedge clk);
#1;data_in = testData5[295];
@(posedge clk);
#1;data_in = testData5[296];
@(posedge clk);
#1;data_in = testData5[297];
@(posedge clk);
#1;data_in = testData5[298];
@(posedge clk);
#1;data_in = testData5[299];
@(posedge clk);
#1;data_in = testData5[300];
@(posedge clk);
#1;data_in = testData5[301];
@(posedge clk);
#1;data_in = testData5[302];
@(posedge clk);
#1;data_in = testData5[303];
@(posedge clk);
#1;data_in = testData5[304];
@(posedge clk);
#1;data_in = testData5[305];
@(posedge clk);
#1;data_in = testData5[306];
@(posedge clk);
#1;data_in = testData5[307];
@(posedge clk);
#1;data_in = testData5[308];
@(posedge clk);
#1;data_in = testData5[309];
@(posedge clk);
#1;data_in = testData5[310];
@(posedge clk);
#1;data_in = testData5[311];
@(posedge clk);
#1;data_in = testData5[312];
@(posedge clk);
#1;data_in = testData5[313];
@(posedge clk);
#1;data_in = testData5[314];
@(posedge clk);
#1;data_in = testData5[315];
@(posedge clk);
#1;data_in = testData5[316];
@(posedge clk);
#1;data_in = testData5[317];
@(posedge clk);
#1;data_in = testData5[318];
@(posedge clk);
#1;data_in = testData5[319];
@(posedge clk);
#1;data_in = testData5[320];
@(posedge clk);
#1;data_in = testData5[321];
@(posedge clk);
#1;data_in = testData5[322];
@(posedge clk);
#1;data_in = testData5[323];
@(posedge clk);
#1;data_in = testData5[324];
@(posedge clk);
#1;data_in = testData5[325];
@(posedge clk);
#1;data_in = testData5[326];
@(posedge clk);
#1;data_in = testData5[327];
@(posedge clk);
#1;data_in = testData5[328];
@(posedge clk);
#1;data_in = testData5[329];
@(posedge clk);
#1;data_in = testData5[330];
@(posedge clk);
#1;data_in = testData5[331];
@(posedge clk);
#1;data_in = testData5[332];
@(posedge clk);
#1;data_in = testData5[333];
@(posedge clk);
#1;data_in = testData5[334];
@(posedge clk);
#1;data_in = testData5[335];
@(posedge clk);
#1;data_in = testData5[336];
@(posedge clk);
#1;data_in = testData5[337];
@(posedge clk);
#1;data_in = testData5[338];
@(posedge clk);
#1;data_in = testData5[339];
@(posedge clk);
#1;data_in = testData5[340];
@(posedge clk);
#1;data_in = testData5[341];
@(posedge clk);
#1;data_in = testData5[342];
@(posedge clk);
#1;data_in = testData5[343];
@(posedge clk);
#1;data_in = testData5[344];
@(posedge clk);
#1;data_in = testData5[345];
@(posedge clk);
#1;data_in = testData5[346];
@(posedge clk);
#1;data_in = testData5[347];
@(posedge clk);
#1;data_in = testData5[348];
@(posedge clk);
#1;data_in = testData5[349];
@(posedge clk);
#1;data_in = testData5[350];
@(posedge clk);
#1;data_in = testData5[351];
@(posedge clk);
#1;data_in = testData5[352];
@(posedge clk);
#1;data_in = testData5[353];
@(posedge clk);
#1;data_in = testData5[354];
@(posedge clk);
#1;data_in = testData5[355];
@(posedge clk);
#1;data_in = testData5[356];
@(posedge clk);
#1;data_in = testData5[357];
@(posedge clk);
#1;data_in = testData5[358];
@(posedge clk);
#1;data_in = testData5[359];
@(posedge clk);
#1;data_in = testData5[360];
@(posedge clk);
#1;data_in = testData5[361];
@(posedge clk);
#1;data_in = testData5[362];
@(posedge clk);
#1;data_in = testData5[363];
@(posedge clk);
#1;data_in = testData5[364];
@(posedge clk);
#1;data_in = testData5[365];
@(posedge clk);
#1;data_in = testData5[366];
@(posedge clk);
#1;data_in = testData5[367];
@(posedge clk);
#1;data_in = testData5[368];
@(posedge clk);
#1;data_in = testData5[369];
@(posedge clk);
#1;data_in = testData5[370];
@(posedge clk);
#1;data_in = testData5[371];
@(posedge clk);
#1;data_in = testData5[372];
@(posedge clk);
#1;data_in = testData5[373];
@(posedge clk);
#1;data_in = testData5[374];
@(posedge clk);
#1;data_in = testData5[375];
@(posedge clk);
#1;data_in = testData5[376];
@(posedge clk);
#1;data_in = testData5[377];
@(posedge clk);
#1;data_in = testData5[378];
@(posedge clk);
#1;data_in = testData5[379];
@(posedge clk);
#1;data_in = testData5[380];
@(posedge clk);
#1;data_in = testData5[381];
@(posedge clk);
#1;data_in = testData5[382];
@(posedge clk);
#1;data_in = testData5[383];
@(posedge clk);
#1;data_in = testData5[384];
@(posedge clk);
#1;data_in = testData5[385];
@(posedge clk);
#1;data_in = testData5[386];
@(posedge clk);
#1;data_in = testData5[387];
@(posedge clk);
#1;data_in = testData5[388];
@(posedge clk);
#1;data_in = testData5[389];
@(posedge clk);
#1;data_in = testData5[390];
@(posedge clk);
#1;data_in = testData5[391];
@(posedge clk);
#1;data_in = testData5[392];
@(posedge clk);
#1;data_in = testData5[393];
@(posedge clk);
#1;data_in = testData5[394];
@(posedge clk);
#1;data_in = testData5[395];
@(posedge clk);
#1;data_in = testData5[396];
@(posedge clk);
#1;data_in = testData5[397];
@(posedge clk);
#1;data_in = testData5[398];
@(posedge clk);
#1;data_in = testData5[399];
@(posedge clk);
#1;data_in = testData5[400];
@(posedge clk);
#1;data_in = testData5[401];
@(posedge clk);
#1;data_in = testData5[402];
@(posedge clk);
#1;data_in = testData5[403];
@(posedge clk);
#1;data_in = testData5[404];
@(posedge clk);
#1;data_in = testData5[405];
@(posedge clk);
#1;data_in = testData5[406];
@(posedge clk);
#1;data_in = testData5[407];
@(posedge clk);
#1;data_in = testData5[408];
@(posedge clk);
#1;data_in = testData5[409];
@(posedge clk);
#1;data_in = testData5[410];
@(posedge clk);
#1;data_in = testData5[411];
@(posedge clk);
#1;data_in = testData5[412];
@(posedge clk);
#1;data_in = testData5[413];
@(posedge clk);
#1;data_in = testData5[414];
@(posedge clk);
#1;data_in = testData5[415];
@(posedge clk);
#1;data_in = testData5[416];
@(posedge clk);
#1;data_in = testData5[417];
@(posedge clk);
#1;data_in = testData5[418];
@(posedge clk);
#1;data_in = testData5[419];
@(posedge clk);
#1;data_in = testData5[420];
@(posedge clk);
#1;data_in = testData5[421];
@(posedge clk);
#1;data_in = testData5[422];
@(posedge clk);
#1;data_in = testData5[423];
@(posedge clk);
#1;data_in = testData5[424];
@(posedge clk);
#1;data_in = testData5[425];
@(posedge clk);
#1;data_in = testData5[426];
@(posedge clk);
#1;data_in = testData5[427];
@(posedge clk);
#1;data_in = testData5[428];
@(posedge clk);
#1;data_in = testData5[429];
@(posedge clk);
#1;data_in = testData5[430];
@(posedge clk);
#1;data_in = testData5[431];
@(posedge clk);
#1;data_in = testData5[432];
@(posedge clk);
#1;data_in = testData5[433];
@(posedge clk);
#1;data_in = testData5[434];
@(posedge clk);
#1;data_in = testData5[435];
@(posedge clk);
#1;data_in = testData5[436];
@(posedge clk);
#1;data_in = testData5[437];
@(posedge clk);
#1;data_in = testData5[438];
@(posedge clk);
#1;data_in = testData5[439];
@(posedge clk);
#1;data_in = testData5[440];
@(posedge clk);
#1;data_in = testData5[441];
@(posedge clk);
#1;data_in = testData5[442];
@(posedge clk);
#1;data_in = testData5[443];
@(posedge clk);
#1;data_in = testData5[444];
@(posedge clk);
#1;data_in = testData5[445];
@(posedge clk);
#1;data_in = testData5[446];
@(posedge clk);
#1;data_in = testData5[447];
@(posedge clk);
#1;data_in = testData5[448];
@(posedge clk);
#1;data_in = testData5[449];
@(posedge clk);
#1;data_in = testData5[450];
@(posedge clk);
#1;data_in = testData5[451];
@(posedge clk);
#1;data_in = testData5[452];
@(posedge clk);
#1;data_in = testData5[453];
@(posedge clk);
#1;data_in = testData5[454];
@(posedge clk);
#1;data_in = testData5[455];
@(posedge clk);
#1;data_in = testData5[456];
@(posedge clk);
#1;data_in = testData5[457];
@(posedge clk);
#1;data_in = testData5[458];
@(posedge clk);
#1;data_in = testData5[459];
@(posedge clk);
#1;data_in = testData5[460];
@(posedge clk);
#1;data_in = testData5[461];
@(posedge clk);
#1;data_in = testData5[462];
@(posedge clk);
#1;data_in = testData5[463];
@(posedge clk);
#1;data_in = testData5[464];
@(posedge clk);
#1;data_in = testData5[465];
@(posedge clk);
#1;data_in = testData5[466];
@(posedge clk);
#1;data_in = testData5[467];
@(posedge clk);
#1;data_in = testData5[468];
@(posedge clk);
#1;data_in = testData5[469];
@(posedge clk);
#1;data_in = testData5[470];
@(posedge clk);
#1;data_in = testData5[471];
@(posedge clk);
#1;data_in = testData5[472];
@(posedge clk);
#1;data_in = testData5[473];
@(posedge clk);
#1;data_in = testData5[474];
@(posedge clk);
#1;data_in = testData5[475];
@(posedge clk);
#1;data_in = testData5[476];
@(posedge clk);
#1;data_in = testData5[477];
@(posedge clk);
#1;data_in = testData5[478];
@(posedge clk);
#1;data_in = testData5[479];
@(posedge clk);
#1;data_in = testData5[480];
@(posedge clk);
#1;data_in = testData5[481];
@(posedge clk);
#1;data_in = testData5[482];
@(posedge clk);
#1;data_in = testData5[483];
@(posedge clk);
#1;data_in = testData5[484];
@(posedge clk);
#1;data_in = testData5[485];
@(posedge clk);
#1;data_in = testData5[486];
@(posedge clk);
#1;data_in = testData5[487];
@(posedge clk);
#1;data_in = testData5[488];
@(posedge clk);
#1;data_in = testData5[489];
@(posedge clk);
#1;data_in = testData5[490];
@(posedge clk);
#1;data_in = testData5[491];
@(posedge clk);
#1;data_in = testData5[492];
@(posedge clk);
#1;data_in = testData5[493];
@(posedge clk);
#1;data_in = testData5[494];
@(posedge clk);
#1;data_in = testData5[495];
@(posedge clk);
#1;data_in = testData5[496];
@(posedge clk);
#1;data_in = testData5[497];
@(posedge clk);
#1;data_in = testData5[498];
@(posedge clk);
#1;data_in = testData5[499];
@(posedge clk);
#1;data_in = testData5[500];
@(posedge clk);
#1;data_in = testData5[501];
@(posedge clk);
#1;data_in = testData5[502];
@(posedge clk);
#1;data_in = testData5[503];
@(posedge clk);
#1;data_in = testData5[504];
@(posedge clk);
#1;data_in = testData5[505];
@(posedge clk);
#1;data_in = testData5[506];
@(posedge clk);
#1;data_in = testData5[507];
@(posedge clk);
#1;data_in = testData5[508];
@(posedge clk);
#1;data_in = testData5[509];
@(posedge clk);
#1;data_in = testData5[510];
@(posedge clk);
#1;data_in = testData5[511];
@(posedge clk);
#1;data_in = testData5[512];
@(posedge clk);
#1;data_in = testData5[513];
@(posedge clk);
#1;data_in = testData5[514];
@(posedge clk);
#1;data_in = testData5[515];
@(posedge clk);
#1;data_in = testData5[516];
@(posedge clk);
#1;data_in = testData5[517];
@(posedge clk);
#1;data_in = testData5[518];
@(posedge clk);
#1;data_in = testData5[519];
@(posedge clk);
#1;data_in = testData5[520];
@(posedge clk);
#1;data_in = testData5[521];
@(posedge clk);
#1;data_in = testData5[522];
@(posedge clk);
#1;data_in = testData5[523];
@(posedge clk);
#1;data_in = testData5[524];
@(posedge clk);
#1;data_in = testData5[525];
@(posedge clk);
#1;data_in = testData5[526];
@(posedge clk);
#1;data_in = testData5[527];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[528]; 
@(posedge clk);
#1;data_in = testData5[529];
@(posedge clk);
#1;data_in = testData5[530];
@(posedge clk);
#1;data_in = testData5[531];
@(posedge clk);
#1;data_in = testData5[532];
@(posedge clk);
#1;data_in = testData5[533];
@(posedge clk);
#1;data_in = testData5[534];
@(posedge clk);
#1;data_in = testData5[535];
@(posedge clk);
#1;data_in = testData5[536];
@(posedge clk);
#1;data_in = testData5[537];
@(posedge clk);
#1;data_in = testData5[538];
@(posedge clk);
#1;data_in = testData5[539];
@(posedge clk);
#1;data_in = testData5[540];
@(posedge clk);
#1;data_in = testData5[541];
@(posedge clk);
#1;data_in = testData5[542];
@(posedge clk);
#1;data_in = testData5[543];
@(posedge clk);
#1;data_in = testData5[544];
@(posedge clk);
#1;data_in = testData5[545];
@(posedge clk);
#1;data_in = testData5[546];
@(posedge clk);
#1;data_in = testData5[547];
@(posedge clk);
#1;data_in = testData5[548];
@(posedge clk);
#1;data_in = testData5[549];
@(posedge clk);
#1;data_in = testData5[550];
@(posedge clk);
#1;data_in = testData5[551];
@(posedge clk);
#1;data_in = testData5[552];
@(posedge clk);
#1;data_in = testData5[553];
@(posedge clk);
#1;data_in = testData5[554];
@(posedge clk);
#1;data_in = testData5[555];
@(posedge clk);
#1;data_in = testData5[556];
@(posedge clk);
#1;data_in = testData5[557];
@(posedge clk);
#1;data_in = testData5[558];
@(posedge clk);
#1;data_in = testData5[559];
@(posedge clk);
#1;data_in = testData5[560];
@(posedge clk);
#1;data_in = testData5[561];
@(posedge clk);
#1;data_in = testData5[562];
@(posedge clk);
#1;data_in = testData5[563];
@(posedge clk);
#1;data_in = testData5[564];
@(posedge clk);
#1;data_in = testData5[565];
@(posedge clk);
#1;data_in = testData5[566];
@(posedge clk);
#1;data_in = testData5[567];
@(posedge clk);
#1;data_in = testData5[568];
@(posedge clk);
#1;data_in = testData5[569];
@(posedge clk);
#1;data_in = testData5[570];
@(posedge clk);
#1;data_in = testData5[571];
@(posedge clk);
#1;data_in = testData5[572];
@(posedge clk);
#1;data_in = testData5[573];
@(posedge clk);
#1;data_in = testData5[574];
@(posedge clk);
#1;data_in = testData5[575];
@(posedge clk);
#1;data_in = testData5[576];
@(posedge clk);
#1;data_in = testData5[577];
@(posedge clk);
#1;data_in = testData5[578];
@(posedge clk);
#1;data_in = testData5[579];
@(posedge clk);
#1;data_in = testData5[580];
@(posedge clk);
#1;data_in = testData5[581];
@(posedge clk);
#1;data_in = testData5[582];
@(posedge clk);
#1;data_in = testData5[583];
@(posedge clk);
#1;data_in = testData5[584];
@(posedge clk);
#1;data_in = testData5[585];
@(posedge clk);
#1;data_in = testData5[586];
@(posedge clk);
#1;data_in = testData5[587];
@(posedge clk);
#1;data_in = testData5[588];
@(posedge clk);
#1;data_in = testData5[589];
@(posedge clk);
#1;data_in = testData5[590];
@(posedge clk);
#1;data_in = testData5[591];
@(posedge clk);
#1;data_in = testData5[592];
@(posedge clk);
#1;data_in = testData5[593];
@(posedge clk);
#1;data_in = testData5[594];
@(posedge clk);
#1;data_in = testData5[595];
@(posedge clk);
#1;data_in = testData5[596];
@(posedge clk);
#1;data_in = testData5[597];
@(posedge clk);
#1;data_in = testData5[598];
@(posedge clk);
#1;data_in = testData5[599];
@(posedge clk);
#1;data_in = testData5[600];
@(posedge clk);
#1;data_in = testData5[601];
@(posedge clk);
#1;data_in = testData5[602];
@(posedge clk);
#1;data_in = testData5[603];
@(posedge clk);
#1;data_in = testData5[604];
@(posedge clk);
#1;data_in = testData5[605];
@(posedge clk);
#1;data_in = testData5[606];
@(posedge clk);
#1;data_in = testData5[607];
@(posedge clk);
#1;data_in = testData5[608];
@(posedge clk);
#1;data_in = testData5[609];
@(posedge clk);
#1;data_in = testData5[610];
@(posedge clk);
#1;data_in = testData5[611];
@(posedge clk);
#1;data_in = testData5[612];
@(posedge clk);
#1;data_in = testData5[613];
@(posedge clk);
#1;data_in = testData5[614];
@(posedge clk);
#1;data_in = testData5[615];
@(posedge clk);
#1;data_in = testData5[616];
@(posedge clk);
#1;data_in = testData5[617];
@(posedge clk);
#1;data_in = testData5[618];
@(posedge clk);
#1;data_in = testData5[619];
@(posedge clk);
#1;data_in = testData5[620];
@(posedge clk);
#1;data_in = testData5[621];
@(posedge clk);
#1;data_in = testData5[622];
@(posedge clk);
#1;data_in = testData5[623];
@(posedge clk);
#1;data_in = testData5[624];
@(posedge clk);
#1;data_in = testData5[625];
@(posedge clk);
#1;data_in = testData5[626];
@(posedge clk);
#1;data_in = testData5[627];
@(posedge clk);
#1;data_in = testData5[628];
@(posedge clk);
#1;data_in = testData5[629];
@(posedge clk);
#1;data_in = testData5[630];
@(posedge clk);
#1;data_in = testData5[631];
@(posedge clk);
#1;data_in = testData5[632];
@(posedge clk);
#1;data_in = testData5[633];
@(posedge clk);
#1;data_in = testData5[634];
@(posedge clk);
#1;data_in = testData5[635];
@(posedge clk);
#1;data_in = testData5[636];
@(posedge clk);
#1;data_in = testData5[637];
@(posedge clk);
#1;data_in = testData5[638];
@(posedge clk);
#1;data_in = testData5[639];
@(posedge clk);
#1;data_in = testData5[640];
@(posedge clk);
#1;data_in = testData5[641];
@(posedge clk);
#1;data_in = testData5[642];
@(posedge clk);
#1;data_in = testData5[643];
@(posedge clk);
#1;data_in = testData5[644];
@(posedge clk);
#1;data_in = testData5[645];
@(posedge clk);
#1;data_in = testData5[646];
@(posedge clk);
#1;data_in = testData5[647];
@(posedge clk);
#1;data_in = testData5[648];
@(posedge clk);
#1;data_in = testData5[649];
@(posedge clk);
#1;data_in = testData5[650];
@(posedge clk);
#1;data_in = testData5[651];
@(posedge clk);
#1;data_in = testData5[652];
@(posedge clk);
#1;data_in = testData5[653];
@(posedge clk);
#1;data_in = testData5[654];
@(posedge clk);
#1;data_in = testData5[655];
@(posedge clk);
#1;data_in = testData5[656];
@(posedge clk);
#1;data_in = testData5[657];
@(posedge clk);
#1;data_in = testData5[658];
@(posedge clk);
#1;data_in = testData5[659];
@(posedge clk);
#1;data_in = testData5[660];
@(posedge clk);
#1;data_in = testData5[661];
@(posedge clk);
#1;data_in = testData5[662];
@(posedge clk);
#1;data_in = testData5[663];
@(posedge clk);
#1;data_in = testData5[664];
@(posedge clk);
#1;data_in = testData5[665];
@(posedge clk);
#1;data_in = testData5[666];
@(posedge clk);
#1;data_in = testData5[667];
@(posedge clk);
#1;data_in = testData5[668];
@(posedge clk);
#1;data_in = testData5[669];
@(posedge clk);
#1;data_in = testData5[670];
@(posedge clk);
#1;data_in = testData5[671];
@(posedge clk);
#1;data_in = testData5[672];
@(posedge clk);
#1;data_in = testData5[673];
@(posedge clk);
#1;data_in = testData5[674];
@(posedge clk);
#1;data_in = testData5[675];
@(posedge clk);
#1;data_in = testData5[676];
@(posedge clk);
#1;data_in = testData5[677];
@(posedge clk);
#1;data_in = testData5[678];
@(posedge clk);
#1;data_in = testData5[679];
@(posedge clk);
#1;data_in = testData5[680];
@(posedge clk);
#1;data_in = testData5[681];
@(posedge clk);
#1;data_in = testData5[682];
@(posedge clk);
#1;data_in = testData5[683];
@(posedge clk);
#1;data_in = testData5[684];
@(posedge clk);
#1;data_in = testData5[685];
@(posedge clk);
#1;data_in = testData5[686];
@(posedge clk);
#1;data_in = testData5[687];
@(posedge clk);
#1;data_in = testData5[688];
@(posedge clk);
#1;data_in = testData5[689];
@(posedge clk);
#1;data_in = testData5[690];
@(posedge clk);
#1;data_in = testData5[691];
@(posedge clk);
#1;data_in = testData5[692];
@(posedge clk);
#1;data_in = testData5[693];
@(posedge clk);
#1;data_in = testData5[694];
@(posedge clk);
#1;data_in = testData5[695];
@(posedge clk);
#1;data_in = testData5[696];
@(posedge clk);
#1;data_in = testData5[697];
@(posedge clk);
#1;data_in = testData5[698];
@(posedge clk);
#1;data_in = testData5[699];
@(posedge clk);
#1;data_in = testData5[700];
@(posedge clk);
#1;data_in = testData5[701];
@(posedge clk);
#1;data_in = testData5[702];
@(posedge clk);
#1;data_in = testData5[703];
@(posedge clk);
#1;data_in = testData5[704];
@(posedge clk);
#1;data_in = testData5[705];
@(posedge clk);
#1;data_in = testData5[706];
@(posedge clk);
#1;data_in = testData5[707];
@(posedge clk);
#1;data_in = testData5[708];
@(posedge clk);
#1;data_in = testData5[709];
@(posedge clk);
#1;data_in = testData5[710];
@(posedge clk);
#1;data_in = testData5[711];
@(posedge clk);
#1;data_in = testData5[712];
@(posedge clk);
#1;data_in = testData5[713];
@(posedge clk);
#1;data_in = testData5[714];
@(posedge clk);
#1;data_in = testData5[715];
@(posedge clk);
#1;data_in = testData5[716];
@(posedge clk);
#1;data_in = testData5[717];
@(posedge clk);
#1;data_in = testData5[718];
@(posedge clk);
#1;data_in = testData5[719];
@(posedge clk);
#1;data_in = testData5[720];
@(posedge clk);
#1;data_in = testData5[721];
@(posedge clk);
#1;data_in = testData5[722];
@(posedge clk);
#1;data_in = testData5[723];
@(posedge clk);
#1;data_in = testData5[724];
@(posedge clk);
#1;data_in = testData5[725];
@(posedge clk);
#1;data_in = testData5[726];
@(posedge clk);
#1;data_in = testData5[727];
@(posedge clk);
#1;data_in = testData5[728];
@(posedge clk);
#1;data_in = testData5[729];
@(posedge clk);
#1;data_in = testData5[730];
@(posedge clk);
#1;data_in = testData5[731];
@(posedge clk);
#1;data_in = testData5[732];
@(posedge clk);
#1;data_in = testData5[733];
@(posedge clk);
#1;data_in = testData5[734];
@(posedge clk);
#1;data_in = testData5[735];
@(posedge clk);
#1;data_in = testData5[736];
@(posedge clk);
#1;data_in = testData5[737];
@(posedge clk);
#1;data_in = testData5[738];
@(posedge clk);
#1;data_in = testData5[739];
@(posedge clk);
#1;data_in = testData5[740];
@(posedge clk);
#1;data_in = testData5[741];
@(posedge clk);
#1;data_in = testData5[742];
@(posedge clk);
#1;data_in = testData5[743];
@(posedge clk);
#1;data_in = testData5[744];
@(posedge clk);
#1;data_in = testData5[745];
@(posedge clk);
#1;data_in = testData5[746];
@(posedge clk);
#1;data_in = testData5[747];
@(posedge clk);
#1;data_in = testData5[748];
@(posedge clk);
#1;data_in = testData5[749];
@(posedge clk);
#1;data_in = testData5[750];
@(posedge clk);
#1;data_in = testData5[751];
@(posedge clk);
#1;data_in = testData5[752];
@(posedge clk);
#1;data_in = testData5[753];
@(posedge clk);
#1;data_in = testData5[754];
@(posedge clk);
#1;data_in = testData5[755];
@(posedge clk);
#1;data_in = testData5[756];
@(posedge clk);
#1;data_in = testData5[757];
@(posedge clk);
#1;data_in = testData5[758];
@(posedge clk);
#1;data_in = testData5[759];
@(posedge clk);
#1;data_in = testData5[760];
@(posedge clk);
#1;data_in = testData5[761];
@(posedge clk);
#1;data_in = testData5[762];
@(posedge clk);
#1;data_in = testData5[763];
@(posedge clk);
#1;data_in = testData5[764];
@(posedge clk);
#1;data_in = testData5[765];
@(posedge clk);
#1;data_in = testData5[766];
@(posedge clk);
#1;data_in = testData5[767];
@(posedge clk);
#1;data_in = testData5[768];
@(posedge clk);
#1;data_in = testData5[769];
@(posedge clk);
#1;data_in = testData5[770];
@(posedge clk);
#1;data_in = testData5[771];
@(posedge clk);
#1;data_in = testData5[772];
@(posedge clk);
#1;data_in = testData5[773];
@(posedge clk);
#1;data_in = testData5[774];
@(posedge clk);
#1;data_in = testData5[775];
@(posedge clk);
#1;data_in = testData5[776];
@(posedge clk);
#1;data_in = testData5[777];
@(posedge clk);
#1;data_in = testData5[778];
@(posedge clk);
#1;data_in = testData5[779];
@(posedge clk);
#1;data_in = testData5[780];
@(posedge clk);
#1;data_in = testData5[781];
@(posedge clk);
#1;data_in = testData5[782];
@(posedge clk);
#1;data_in = testData5[783];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[784]; 
@(posedge clk);
#1;data_in = testData5[785];
@(posedge clk);
#1;data_in = testData5[786];
@(posedge clk);
#1;data_in = testData5[787];
@(posedge clk);
#1;data_in = testData5[788];
@(posedge clk);
#1;data_in = testData5[789];
@(posedge clk);
#1;data_in = testData5[790];
@(posedge clk);
#1;data_in = testData5[791];
@(posedge clk);
#1;data_in = testData5[792];
@(posedge clk);
#1;data_in = testData5[793];
@(posedge clk);
#1;data_in = testData5[794];
@(posedge clk);
#1;data_in = testData5[795];
@(posedge clk);
#1;data_in = testData5[796];
@(posedge clk);
#1;data_in = testData5[797];
@(posedge clk);
#1;data_in = testData5[798];
@(posedge clk);
#1;data_in = testData5[799];
@(posedge clk);
#1;data_in = testData5[800];
@(posedge clk);
#1;data_in = testData5[801];
@(posedge clk);
#1;data_in = testData5[802];
@(posedge clk);
#1;data_in = testData5[803];
@(posedge clk);
#1;data_in = testData5[804];
@(posedge clk);
#1;data_in = testData5[805];
@(posedge clk);
#1;data_in = testData5[806];
@(posedge clk);
#1;data_in = testData5[807];
@(posedge clk);
#1;data_in = testData5[808];
@(posedge clk);
#1;data_in = testData5[809];
@(posedge clk);
#1;data_in = testData5[810];
@(posedge clk);
#1;data_in = testData5[811];
@(posedge clk);
#1;data_in = testData5[812];
@(posedge clk);
#1;data_in = testData5[813];
@(posedge clk);
#1;data_in = testData5[814];
@(posedge clk);
#1;data_in = testData5[815];
@(posedge clk);
#1;data_in = testData5[816];
@(posedge clk);
#1;data_in = testData5[817];
@(posedge clk);
#1;data_in = testData5[818];
@(posedge clk);
#1;data_in = testData5[819];
@(posedge clk);
#1;data_in = testData5[820];
@(posedge clk);
#1;data_in = testData5[821];
@(posedge clk);
#1;data_in = testData5[822];
@(posedge clk);
#1;data_in = testData5[823];
@(posedge clk);
#1;data_in = testData5[824];
@(posedge clk);
#1;data_in = testData5[825];
@(posedge clk);
#1;data_in = testData5[826];
@(posedge clk);
#1;data_in = testData5[827];
@(posedge clk);
#1;data_in = testData5[828];
@(posedge clk);
#1;data_in = testData5[829];
@(posedge clk);
#1;data_in = testData5[830];
@(posedge clk);
#1;data_in = testData5[831];
@(posedge clk);
#1;data_in = testData5[832];
@(posedge clk);
#1;data_in = testData5[833];
@(posedge clk);
#1;data_in = testData5[834];
@(posedge clk);
#1;data_in = testData5[835];
@(posedge clk);
#1;data_in = testData5[836];
@(posedge clk);
#1;data_in = testData5[837];
@(posedge clk);
#1;data_in = testData5[838];
@(posedge clk);
#1;data_in = testData5[839];
@(posedge clk);
#1;data_in = testData5[840];
@(posedge clk);
#1;data_in = testData5[841];
@(posedge clk);
#1;data_in = testData5[842];
@(posedge clk);
#1;data_in = testData5[843];
@(posedge clk);
#1;data_in = testData5[844];
@(posedge clk);
#1;data_in = testData5[845];
@(posedge clk);
#1;data_in = testData5[846];
@(posedge clk);
#1;data_in = testData5[847];
@(posedge clk);
#1;data_in = testData5[848];
@(posedge clk);
#1;data_in = testData5[849];
@(posedge clk);
#1;data_in = testData5[850];
@(posedge clk);
#1;data_in = testData5[851];
@(posedge clk);
#1;data_in = testData5[852];
@(posedge clk);
#1;data_in = testData5[853];
@(posedge clk);
#1;data_in = testData5[854];
@(posedge clk);
#1;data_in = testData5[855];
@(posedge clk);
#1;data_in = testData5[856];
@(posedge clk);
#1;data_in = testData5[857];
@(posedge clk);
#1;data_in = testData5[858];
@(posedge clk);
#1;data_in = testData5[859];
@(posedge clk);
#1;data_in = testData5[860];
@(posedge clk);
#1;data_in = testData5[861];
@(posedge clk);
#1;data_in = testData5[862];
@(posedge clk);
#1;data_in = testData5[863];
@(posedge clk);
#1;data_in = testData5[864];
@(posedge clk);
#1;data_in = testData5[865];
@(posedge clk);
#1;data_in = testData5[866];
@(posedge clk);
#1;data_in = testData5[867];
@(posedge clk);
#1;data_in = testData5[868];
@(posedge clk);
#1;data_in = testData5[869];
@(posedge clk);
#1;data_in = testData5[870];
@(posedge clk);
#1;data_in = testData5[871];
@(posedge clk);
#1;data_in = testData5[872];
@(posedge clk);
#1;data_in = testData5[873];
@(posedge clk);
#1;data_in = testData5[874];
@(posedge clk);
#1;data_in = testData5[875];
@(posedge clk);
#1;data_in = testData5[876];
@(posedge clk);
#1;data_in = testData5[877];
@(posedge clk);
#1;data_in = testData5[878];
@(posedge clk);
#1;data_in = testData5[879];
@(posedge clk);
#1;data_in = testData5[880];
@(posedge clk);
#1;data_in = testData5[881];
@(posedge clk);
#1;data_in = testData5[882];
@(posedge clk);
#1;data_in = testData5[883];
@(posedge clk);
#1;data_in = testData5[884];
@(posedge clk);
#1;data_in = testData5[885];
@(posedge clk);
#1;data_in = testData5[886];
@(posedge clk);
#1;data_in = testData5[887];
@(posedge clk);
#1;data_in = testData5[888];
@(posedge clk);
#1;data_in = testData5[889];
@(posedge clk);
#1;data_in = testData5[890];
@(posedge clk);
#1;data_in = testData5[891];
@(posedge clk);
#1;data_in = testData5[892];
@(posedge clk);
#1;data_in = testData5[893];
@(posedge clk);
#1;data_in = testData5[894];
@(posedge clk);
#1;data_in = testData5[895];
@(posedge clk);
#1;data_in = testData5[896];
@(posedge clk);
#1;data_in = testData5[897];
@(posedge clk);
#1;data_in = testData5[898];
@(posedge clk);
#1;data_in = testData5[899];
@(posedge clk);
#1;data_in = testData5[900];
@(posedge clk);
#1;data_in = testData5[901];
@(posedge clk);
#1;data_in = testData5[902];
@(posedge clk);
#1;data_in = testData5[903];
@(posedge clk);
#1;data_in = testData5[904];
@(posedge clk);
#1;data_in = testData5[905];
@(posedge clk);
#1;data_in = testData5[906];
@(posedge clk);
#1;data_in = testData5[907];
@(posedge clk);
#1;data_in = testData5[908];
@(posedge clk);
#1;data_in = testData5[909];
@(posedge clk);
#1;data_in = testData5[910];
@(posedge clk);
#1;data_in = testData5[911];
@(posedge clk);
#1;data_in = testData5[912];
@(posedge clk);
#1;data_in = testData5[913];
@(posedge clk);
#1;data_in = testData5[914];
@(posedge clk);
#1;data_in = testData5[915];
@(posedge clk);
#1;data_in = testData5[916];
@(posedge clk);
#1;data_in = testData5[917];
@(posedge clk);
#1;data_in = testData5[918];
@(posedge clk);
#1;data_in = testData5[919];
@(posedge clk);
#1;data_in = testData5[920];
@(posedge clk);
#1;data_in = testData5[921];
@(posedge clk);
#1;data_in = testData5[922];
@(posedge clk);
#1;data_in = testData5[923];
@(posedge clk);
#1;data_in = testData5[924];
@(posedge clk);
#1;data_in = testData5[925];
@(posedge clk);
#1;data_in = testData5[926];
@(posedge clk);
#1;data_in = testData5[927];
@(posedge clk);
#1;data_in = testData5[928];
@(posedge clk);
#1;data_in = testData5[929];
@(posedge clk);
#1;data_in = testData5[930];
@(posedge clk);
#1;data_in = testData5[931];
@(posedge clk);
#1;data_in = testData5[932];
@(posedge clk);
#1;data_in = testData5[933];
@(posedge clk);
#1;data_in = testData5[934];
@(posedge clk);
#1;data_in = testData5[935];
@(posedge clk);
#1;data_in = testData5[936];
@(posedge clk);
#1;data_in = testData5[937];
@(posedge clk);
#1;data_in = testData5[938];
@(posedge clk);
#1;data_in = testData5[939];
@(posedge clk);
#1;data_in = testData5[940];
@(posedge clk);
#1;data_in = testData5[941];
@(posedge clk);
#1;data_in = testData5[942];
@(posedge clk);
#1;data_in = testData5[943];
@(posedge clk);
#1;data_in = testData5[944];
@(posedge clk);
#1;data_in = testData5[945];
@(posedge clk);
#1;data_in = testData5[946];
@(posedge clk);
#1;data_in = testData5[947];
@(posedge clk);
#1;data_in = testData5[948];
@(posedge clk);
#1;data_in = testData5[949];
@(posedge clk);
#1;data_in = testData5[950];
@(posedge clk);
#1;data_in = testData5[951];
@(posedge clk);
#1;data_in = testData5[952];
@(posedge clk);
#1;data_in = testData5[953];
@(posedge clk);
#1;data_in = testData5[954];
@(posedge clk);
#1;data_in = testData5[955];
@(posedge clk);
#1;data_in = testData5[956];
@(posedge clk);
#1;data_in = testData5[957];
@(posedge clk);
#1;data_in = testData5[958];
@(posedge clk);
#1;data_in = testData5[959];
@(posedge clk);
#1;data_in = testData5[960];
@(posedge clk);
#1;data_in = testData5[961];
@(posedge clk);
#1;data_in = testData5[962];
@(posedge clk);
#1;data_in = testData5[963];
@(posedge clk);
#1;data_in = testData5[964];
@(posedge clk);
#1;data_in = testData5[965];
@(posedge clk);
#1;data_in = testData5[966];
@(posedge clk);
#1;data_in = testData5[967];
@(posedge clk);
#1;data_in = testData5[968];
@(posedge clk);
#1;data_in = testData5[969];
@(posedge clk);
#1;data_in = testData5[970];
@(posedge clk);
#1;data_in = testData5[971];
@(posedge clk);
#1;data_in = testData5[972];
@(posedge clk);
#1;data_in = testData5[973];
@(posedge clk);
#1;data_in = testData5[974];
@(posedge clk);
#1;data_in = testData5[975];
@(posedge clk);
#1;data_in = testData5[976];
@(posedge clk);
#1;data_in = testData5[977];
@(posedge clk);
#1;data_in = testData5[978];
@(posedge clk);
#1;data_in = testData5[979];
@(posedge clk);
#1;data_in = testData5[980];
@(posedge clk);
#1;data_in = testData5[981];
@(posedge clk);
#1;data_in = testData5[982];
@(posedge clk);
#1;data_in = testData5[983];
@(posedge clk);
#1;data_in = testData5[984];
@(posedge clk);
#1;data_in = testData5[985];
@(posedge clk);
#1;data_in = testData5[986];
@(posedge clk);
#1;data_in = testData5[987];
@(posedge clk);
#1;data_in = testData5[988];
@(posedge clk);
#1;data_in = testData5[989];
@(posedge clk);
#1;data_in = testData5[990];
@(posedge clk);
#1;data_in = testData5[991];
@(posedge clk);
#1;data_in = testData5[992];
@(posedge clk);
#1;data_in = testData5[993];
@(posedge clk);
#1;data_in = testData5[994];
@(posedge clk);
#1;data_in = testData5[995];
@(posedge clk);
#1;data_in = testData5[996];
@(posedge clk);
#1;data_in = testData5[997];
@(posedge clk);
#1;data_in = testData5[998];
@(posedge clk);
#1;data_in = testData5[999];
@(posedge clk);
#1;data_in = testData5[1000];
@(posedge clk);
#1;data_in = testData5[1001];
@(posedge clk);
#1;data_in = testData5[1002];
@(posedge clk);
#1;data_in = testData5[1003];
@(posedge clk);
#1;data_in = testData5[1004];
@(posedge clk);
#1;data_in = testData5[1005];
@(posedge clk);
#1;data_in = testData5[1006];
@(posedge clk);
#1;data_in = testData5[1007];
@(posedge clk);
#1;data_in = testData5[1008];
@(posedge clk);
#1;data_in = testData5[1009];
@(posedge clk);
#1;data_in = testData5[1010];
@(posedge clk);
#1;data_in = testData5[1011];
@(posedge clk);
#1;data_in = testData5[1012];
@(posedge clk);
#1;data_in = testData5[1013];
@(posedge clk);
#1;data_in = testData5[1014];
@(posedge clk);
#1;data_in = testData5[1015];
@(posedge clk);
#1;data_in = testData5[1016];
@(posedge clk);
#1;data_in = testData5[1017];
@(posedge clk);
#1;data_in = testData5[1018];
@(posedge clk);
#1;data_in = testData5[1019];
@(posedge clk);
#1;data_in = testData5[1020];
@(posedge clk);
#1;data_in = testData5[1021];
@(posedge clk);
#1;data_in = testData5[1022];
@(posedge clk);
#1;data_in = testData5[1023];
@(posedge clk);
#1;data_in = testData5[1024];
@(posedge clk);
#1;data_in = testData5[1025];
@(posedge clk);
#1;data_in = testData5[1026];
@(posedge clk);
#1;data_in = testData5[1027];
@(posedge clk);
#1;data_in = testData5[1028];
@(posedge clk);
#1;data_in = testData5[1029];
@(posedge clk);
#1;data_in = testData5[1030];
@(posedge clk);
#1;data_in = testData5[1031];
@(posedge clk);
#1;data_in = testData5[1032];
@(posedge clk);
#1;data_in = testData5[1033];
@(posedge clk);
#1;data_in = testData5[1034];
@(posedge clk);
#1;data_in = testData5[1035];
@(posedge clk);
#1;data_in = testData5[1036];
@(posedge clk);
#1;data_in = testData5[1037];
@(posedge clk);
#1;data_in = testData5[1038];
@(posedge clk);
#1;data_in = testData5[1039];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1040]; 
@(posedge clk);
#1;data_in = testData5[1041];
@(posedge clk);
#1;data_in = testData5[1042];
@(posedge clk);
#1;data_in = testData5[1043];
@(posedge clk);
#1;data_in = testData5[1044];
@(posedge clk);
#1;data_in = testData5[1045];
@(posedge clk);
#1;data_in = testData5[1046];
@(posedge clk);
#1;data_in = testData5[1047];
@(posedge clk);
#1;data_in = testData5[1048];
@(posedge clk);
#1;data_in = testData5[1049];
@(posedge clk);
#1;data_in = testData5[1050];
@(posedge clk);
#1;data_in = testData5[1051];
@(posedge clk);
#1;data_in = testData5[1052];
@(posedge clk);
#1;data_in = testData5[1053];
@(posedge clk);
#1;data_in = testData5[1054];
@(posedge clk);
#1;data_in = testData5[1055];
@(posedge clk);
#1;data_in = testData5[1056];
@(posedge clk);
#1;data_in = testData5[1057];
@(posedge clk);
#1;data_in = testData5[1058];
@(posedge clk);
#1;data_in = testData5[1059];
@(posedge clk);
#1;data_in = testData5[1060];
@(posedge clk);
#1;data_in = testData5[1061];
@(posedge clk);
#1;data_in = testData5[1062];
@(posedge clk);
#1;data_in = testData5[1063];
@(posedge clk);
#1;data_in = testData5[1064];
@(posedge clk);
#1;data_in = testData5[1065];
@(posedge clk);
#1;data_in = testData5[1066];
@(posedge clk);
#1;data_in = testData5[1067];
@(posedge clk);
#1;data_in = testData5[1068];
@(posedge clk);
#1;data_in = testData5[1069];
@(posedge clk);
#1;data_in = testData5[1070];
@(posedge clk);
#1;data_in = testData5[1071];
@(posedge clk);
#1;data_in = testData5[1072];
@(posedge clk);
#1;data_in = testData5[1073];
@(posedge clk);
#1;data_in = testData5[1074];
@(posedge clk);
#1;data_in = testData5[1075];
@(posedge clk);
#1;data_in = testData5[1076];
@(posedge clk);
#1;data_in = testData5[1077];
@(posedge clk);
#1;data_in = testData5[1078];
@(posedge clk);
#1;data_in = testData5[1079];
@(posedge clk);
#1;data_in = testData5[1080];
@(posedge clk);
#1;data_in = testData5[1081];
@(posedge clk);
#1;data_in = testData5[1082];
@(posedge clk);
#1;data_in = testData5[1083];
@(posedge clk);
#1;data_in = testData5[1084];
@(posedge clk);
#1;data_in = testData5[1085];
@(posedge clk);
#1;data_in = testData5[1086];
@(posedge clk);
#1;data_in = testData5[1087];
@(posedge clk);
#1;data_in = testData5[1088];
@(posedge clk);
#1;data_in = testData5[1089];
@(posedge clk);
#1;data_in = testData5[1090];
@(posedge clk);
#1;data_in = testData5[1091];
@(posedge clk);
#1;data_in = testData5[1092];
@(posedge clk);
#1;data_in = testData5[1093];
@(posedge clk);
#1;data_in = testData5[1094];
@(posedge clk);
#1;data_in = testData5[1095];
@(posedge clk);
#1;data_in = testData5[1096];
@(posedge clk);
#1;data_in = testData5[1097];
@(posedge clk);
#1;data_in = testData5[1098];
@(posedge clk);
#1;data_in = testData5[1099];
@(posedge clk);
#1;data_in = testData5[1100];
@(posedge clk);
#1;data_in = testData5[1101];
@(posedge clk);
#1;data_in = testData5[1102];
@(posedge clk);
#1;data_in = testData5[1103];
@(posedge clk);
#1;data_in = testData5[1104];
@(posedge clk);
#1;data_in = testData5[1105];
@(posedge clk);
#1;data_in = testData5[1106];
@(posedge clk);
#1;data_in = testData5[1107];
@(posedge clk);
#1;data_in = testData5[1108];
@(posedge clk);
#1;data_in = testData5[1109];
@(posedge clk);
#1;data_in = testData5[1110];
@(posedge clk);
#1;data_in = testData5[1111];
@(posedge clk);
#1;data_in = testData5[1112];
@(posedge clk);
#1;data_in = testData5[1113];
@(posedge clk);
#1;data_in = testData5[1114];
@(posedge clk);
#1;data_in = testData5[1115];
@(posedge clk);
#1;data_in = testData5[1116];
@(posedge clk);
#1;data_in = testData5[1117];
@(posedge clk);
#1;data_in = testData5[1118];
@(posedge clk);
#1;data_in = testData5[1119];
@(posedge clk);
#1;data_in = testData5[1120];
@(posedge clk);
#1;data_in = testData5[1121];
@(posedge clk);
#1;data_in = testData5[1122];
@(posedge clk);
#1;data_in = testData5[1123];
@(posedge clk);
#1;data_in = testData5[1124];
@(posedge clk);
#1;data_in = testData5[1125];
@(posedge clk);
#1;data_in = testData5[1126];
@(posedge clk);
#1;data_in = testData5[1127];
@(posedge clk);
#1;data_in = testData5[1128];
@(posedge clk);
#1;data_in = testData5[1129];
@(posedge clk);
#1;data_in = testData5[1130];
@(posedge clk);
#1;data_in = testData5[1131];
@(posedge clk);
#1;data_in = testData5[1132];
@(posedge clk);
#1;data_in = testData5[1133];
@(posedge clk);
#1;data_in = testData5[1134];
@(posedge clk);
#1;data_in = testData5[1135];
@(posedge clk);
#1;data_in = testData5[1136];
@(posedge clk);
#1;data_in = testData5[1137];
@(posedge clk);
#1;data_in = testData5[1138];
@(posedge clk);
#1;data_in = testData5[1139];
@(posedge clk);
#1;data_in = testData5[1140];
@(posedge clk);
#1;data_in = testData5[1141];
@(posedge clk);
#1;data_in = testData5[1142];
@(posedge clk);
#1;data_in = testData5[1143];
@(posedge clk);
#1;data_in = testData5[1144];
@(posedge clk);
#1;data_in = testData5[1145];
@(posedge clk);
#1;data_in = testData5[1146];
@(posedge clk);
#1;data_in = testData5[1147];
@(posedge clk);
#1;data_in = testData5[1148];
@(posedge clk);
#1;data_in = testData5[1149];
@(posedge clk);
#1;data_in = testData5[1150];
@(posedge clk);
#1;data_in = testData5[1151];
@(posedge clk);
#1;data_in = testData5[1152];
@(posedge clk);
#1;data_in = testData5[1153];
@(posedge clk);
#1;data_in = testData5[1154];
@(posedge clk);
#1;data_in = testData5[1155];
@(posedge clk);
#1;data_in = testData5[1156];
@(posedge clk);
#1;data_in = testData5[1157];
@(posedge clk);
#1;data_in = testData5[1158];
@(posedge clk);
#1;data_in = testData5[1159];
@(posedge clk);
#1;data_in = testData5[1160];
@(posedge clk);
#1;data_in = testData5[1161];
@(posedge clk);
#1;data_in = testData5[1162];
@(posedge clk);
#1;data_in = testData5[1163];
@(posedge clk);
#1;data_in = testData5[1164];
@(posedge clk);
#1;data_in = testData5[1165];
@(posedge clk);
#1;data_in = testData5[1166];
@(posedge clk);
#1;data_in = testData5[1167];
@(posedge clk);
#1;data_in = testData5[1168];
@(posedge clk);
#1;data_in = testData5[1169];
@(posedge clk);
#1;data_in = testData5[1170];
@(posedge clk);
#1;data_in = testData5[1171];
@(posedge clk);
#1;data_in = testData5[1172];
@(posedge clk);
#1;data_in = testData5[1173];
@(posedge clk);
#1;data_in = testData5[1174];
@(posedge clk);
#1;data_in = testData5[1175];
@(posedge clk);
#1;data_in = testData5[1176];
@(posedge clk);
#1;data_in = testData5[1177];
@(posedge clk);
#1;data_in = testData5[1178];
@(posedge clk);
#1;data_in = testData5[1179];
@(posedge clk);
#1;data_in = testData5[1180];
@(posedge clk);
#1;data_in = testData5[1181];
@(posedge clk);
#1;data_in = testData5[1182];
@(posedge clk);
#1;data_in = testData5[1183];
@(posedge clk);
#1;data_in = testData5[1184];
@(posedge clk);
#1;data_in = testData5[1185];
@(posedge clk);
#1;data_in = testData5[1186];
@(posedge clk);
#1;data_in = testData5[1187];
@(posedge clk);
#1;data_in = testData5[1188];
@(posedge clk);
#1;data_in = testData5[1189];
@(posedge clk);
#1;data_in = testData5[1190];
@(posedge clk);
#1;data_in = testData5[1191];
@(posedge clk);
#1;data_in = testData5[1192];
@(posedge clk);
#1;data_in = testData5[1193];
@(posedge clk);
#1;data_in = testData5[1194];
@(posedge clk);
#1;data_in = testData5[1195];
@(posedge clk);
#1;data_in = testData5[1196];
@(posedge clk);
#1;data_in = testData5[1197];
@(posedge clk);
#1;data_in = testData5[1198];
@(posedge clk);
#1;data_in = testData5[1199];
@(posedge clk);
#1;data_in = testData5[1200];
@(posedge clk);
#1;data_in = testData5[1201];
@(posedge clk);
#1;data_in = testData5[1202];
@(posedge clk);
#1;data_in = testData5[1203];
@(posedge clk);
#1;data_in = testData5[1204];
@(posedge clk);
#1;data_in = testData5[1205];
@(posedge clk);
#1;data_in = testData5[1206];
@(posedge clk);
#1;data_in = testData5[1207];
@(posedge clk);
#1;data_in = testData5[1208];
@(posedge clk);
#1;data_in = testData5[1209];
@(posedge clk);
#1;data_in = testData5[1210];
@(posedge clk);
#1;data_in = testData5[1211];
@(posedge clk);
#1;data_in = testData5[1212];
@(posedge clk);
#1;data_in = testData5[1213];
@(posedge clk);
#1;data_in = testData5[1214];
@(posedge clk);
#1;data_in = testData5[1215];
@(posedge clk);
#1;data_in = testData5[1216];
@(posedge clk);
#1;data_in = testData5[1217];
@(posedge clk);
#1;data_in = testData5[1218];
@(posedge clk);
#1;data_in = testData5[1219];
@(posedge clk);
#1;data_in = testData5[1220];
@(posedge clk);
#1;data_in = testData5[1221];
@(posedge clk);
#1;data_in = testData5[1222];
@(posedge clk);
#1;data_in = testData5[1223];
@(posedge clk);
#1;data_in = testData5[1224];
@(posedge clk);
#1;data_in = testData5[1225];
@(posedge clk);
#1;data_in = testData5[1226];
@(posedge clk);
#1;data_in = testData5[1227];
@(posedge clk);
#1;data_in = testData5[1228];
@(posedge clk);
#1;data_in = testData5[1229];
@(posedge clk);
#1;data_in = testData5[1230];
@(posedge clk);
#1;data_in = testData5[1231];
@(posedge clk);
#1;data_in = testData5[1232];
@(posedge clk);
#1;data_in = testData5[1233];
@(posedge clk);
#1;data_in = testData5[1234];
@(posedge clk);
#1;data_in = testData5[1235];
@(posedge clk);
#1;data_in = testData5[1236];
@(posedge clk);
#1;data_in = testData5[1237];
@(posedge clk);
#1;data_in = testData5[1238];
@(posedge clk);
#1;data_in = testData5[1239];
@(posedge clk);
#1;data_in = testData5[1240];
@(posedge clk);
#1;data_in = testData5[1241];
@(posedge clk);
#1;data_in = testData5[1242];
@(posedge clk);
#1;data_in = testData5[1243];
@(posedge clk);
#1;data_in = testData5[1244];
@(posedge clk);
#1;data_in = testData5[1245];
@(posedge clk);
#1;data_in = testData5[1246];
@(posedge clk);
#1;data_in = testData5[1247];
@(posedge clk);
#1;data_in = testData5[1248];
@(posedge clk);
#1;data_in = testData5[1249];
@(posedge clk);
#1;data_in = testData5[1250];
@(posedge clk);
#1;data_in = testData5[1251];
@(posedge clk);
#1;data_in = testData5[1252];
@(posedge clk);
#1;data_in = testData5[1253];
@(posedge clk);
#1;data_in = testData5[1254];
@(posedge clk);
#1;data_in = testData5[1255];
@(posedge clk);
#1;data_in = testData5[1256];
@(posedge clk);
#1;data_in = testData5[1257];
@(posedge clk);
#1;data_in = testData5[1258];
@(posedge clk);
#1;data_in = testData5[1259];
@(posedge clk);
#1;data_in = testData5[1260];
@(posedge clk);
#1;data_in = testData5[1261];
@(posedge clk);
#1;data_in = testData5[1262];
@(posedge clk);
#1;data_in = testData5[1263];
@(posedge clk);
#1;data_in = testData5[1264];
@(posedge clk);
#1;data_in = testData5[1265];
@(posedge clk);
#1;data_in = testData5[1266];
@(posedge clk);
#1;data_in = testData5[1267];
@(posedge clk);
#1;data_in = testData5[1268];
@(posedge clk);
#1;data_in = testData5[1269];
@(posedge clk);
#1;data_in = testData5[1270];
@(posedge clk);
#1;data_in = testData5[1271];
@(posedge clk);
#1;data_in = testData5[1272];
@(posedge clk);
#1;data_in = testData5[1273];
@(posedge clk);
#1;data_in = testData5[1274];
@(posedge clk);
#1;data_in = testData5[1275];
@(posedge clk);
#1;data_in = testData5[1276];
@(posedge clk);
#1;data_in = testData5[1277];
@(posedge clk);
#1;data_in = testData5[1278];
@(posedge clk);
#1;data_in = testData5[1279];
@(posedge clk);
#1;data_in = testData5[1280];
@(posedge clk);
#1;data_in = testData5[1281];
@(posedge clk);
#1;data_in = testData5[1282];
@(posedge clk);
#1;data_in = testData5[1283];
@(posedge clk);
#1;data_in = testData5[1284];
@(posedge clk);
#1;data_in = testData5[1285];
@(posedge clk);
#1;data_in = testData5[1286];
@(posedge clk);
#1;data_in = testData5[1287];
@(posedge clk);
#1;data_in = testData5[1288];
@(posedge clk);
#1;data_in = testData5[1289];
@(posedge clk);
#1;data_in = testData5[1290];
@(posedge clk);
#1;data_in = testData5[1291];
@(posedge clk);
#1;data_in = testData5[1292];
@(posedge clk);
#1;data_in = testData5[1293];
@(posedge clk);
#1;data_in = testData5[1294];
@(posedge clk);
#1;data_in = testData5[1295];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1296]; 
@(posedge clk);
#1;data_in = testData5[1297];
@(posedge clk);
#1;data_in = testData5[1298];
@(posedge clk);
#1;data_in = testData5[1299];
@(posedge clk);
#1;data_in = testData5[1300];
@(posedge clk);
#1;data_in = testData5[1301];
@(posedge clk);
#1;data_in = testData5[1302];
@(posedge clk);
#1;data_in = testData5[1303];
@(posedge clk);
#1;data_in = testData5[1304];
@(posedge clk);
#1;data_in = testData5[1305];
@(posedge clk);
#1;data_in = testData5[1306];
@(posedge clk);
#1;data_in = testData5[1307];
@(posedge clk);
#1;data_in = testData5[1308];
@(posedge clk);
#1;data_in = testData5[1309];
@(posedge clk);
#1;data_in = testData5[1310];
@(posedge clk);
#1;data_in = testData5[1311];
@(posedge clk);
#1;data_in = testData5[1312];
@(posedge clk);
#1;data_in = testData5[1313];
@(posedge clk);
#1;data_in = testData5[1314];
@(posedge clk);
#1;data_in = testData5[1315];
@(posedge clk);
#1;data_in = testData5[1316];
@(posedge clk);
#1;data_in = testData5[1317];
@(posedge clk);
#1;data_in = testData5[1318];
@(posedge clk);
#1;data_in = testData5[1319];
@(posedge clk);
#1;data_in = testData5[1320];
@(posedge clk);
#1;data_in = testData5[1321];
@(posedge clk);
#1;data_in = testData5[1322];
@(posedge clk);
#1;data_in = testData5[1323];
@(posedge clk);
#1;data_in = testData5[1324];
@(posedge clk);
#1;data_in = testData5[1325];
@(posedge clk);
#1;data_in = testData5[1326];
@(posedge clk);
#1;data_in = testData5[1327];
@(posedge clk);
#1;data_in = testData5[1328];
@(posedge clk);
#1;data_in = testData5[1329];
@(posedge clk);
#1;data_in = testData5[1330];
@(posedge clk);
#1;data_in = testData5[1331];
@(posedge clk);
#1;data_in = testData5[1332];
@(posedge clk);
#1;data_in = testData5[1333];
@(posedge clk);
#1;data_in = testData5[1334];
@(posedge clk);
#1;data_in = testData5[1335];
@(posedge clk);
#1;data_in = testData5[1336];
@(posedge clk);
#1;data_in = testData5[1337];
@(posedge clk);
#1;data_in = testData5[1338];
@(posedge clk);
#1;data_in = testData5[1339];
@(posedge clk);
#1;data_in = testData5[1340];
@(posedge clk);
#1;data_in = testData5[1341];
@(posedge clk);
#1;data_in = testData5[1342];
@(posedge clk);
#1;data_in = testData5[1343];
@(posedge clk);
#1;data_in = testData5[1344];
@(posedge clk);
#1;data_in = testData5[1345];
@(posedge clk);
#1;data_in = testData5[1346];
@(posedge clk);
#1;data_in = testData5[1347];
@(posedge clk);
#1;data_in = testData5[1348];
@(posedge clk);
#1;data_in = testData5[1349];
@(posedge clk);
#1;data_in = testData5[1350];
@(posedge clk);
#1;data_in = testData5[1351];
@(posedge clk);
#1;data_in = testData5[1352];
@(posedge clk);
#1;data_in = testData5[1353];
@(posedge clk);
#1;data_in = testData5[1354];
@(posedge clk);
#1;data_in = testData5[1355];
@(posedge clk);
#1;data_in = testData5[1356];
@(posedge clk);
#1;data_in = testData5[1357];
@(posedge clk);
#1;data_in = testData5[1358];
@(posedge clk);
#1;data_in = testData5[1359];
@(posedge clk);
#1;data_in = testData5[1360];
@(posedge clk);
#1;data_in = testData5[1361];
@(posedge clk);
#1;data_in = testData5[1362];
@(posedge clk);
#1;data_in = testData5[1363];
@(posedge clk);
#1;data_in = testData5[1364];
@(posedge clk);
#1;data_in = testData5[1365];
@(posedge clk);
#1;data_in = testData5[1366];
@(posedge clk);
#1;data_in = testData5[1367];
@(posedge clk);
#1;data_in = testData5[1368];
@(posedge clk);
#1;data_in = testData5[1369];
@(posedge clk);
#1;data_in = testData5[1370];
@(posedge clk);
#1;data_in = testData5[1371];
@(posedge clk);
#1;data_in = testData5[1372];
@(posedge clk);
#1;data_in = testData5[1373];
@(posedge clk);
#1;data_in = testData5[1374];
@(posedge clk);
#1;data_in = testData5[1375];
@(posedge clk);
#1;data_in = testData5[1376];
@(posedge clk);
#1;data_in = testData5[1377];
@(posedge clk);
#1;data_in = testData5[1378];
@(posedge clk);
#1;data_in = testData5[1379];
@(posedge clk);
#1;data_in = testData5[1380];
@(posedge clk);
#1;data_in = testData5[1381];
@(posedge clk);
#1;data_in = testData5[1382];
@(posedge clk);
#1;data_in = testData5[1383];
@(posedge clk);
#1;data_in = testData5[1384];
@(posedge clk);
#1;data_in = testData5[1385];
@(posedge clk);
#1;data_in = testData5[1386];
@(posedge clk);
#1;data_in = testData5[1387];
@(posedge clk);
#1;data_in = testData5[1388];
@(posedge clk);
#1;data_in = testData5[1389];
@(posedge clk);
#1;data_in = testData5[1390];
@(posedge clk);
#1;data_in = testData5[1391];
@(posedge clk);
#1;data_in = testData5[1392];
@(posedge clk);
#1;data_in = testData5[1393];
@(posedge clk);
#1;data_in = testData5[1394];
@(posedge clk);
#1;data_in = testData5[1395];
@(posedge clk);
#1;data_in = testData5[1396];
@(posedge clk);
#1;data_in = testData5[1397];
@(posedge clk);
#1;data_in = testData5[1398];
@(posedge clk);
#1;data_in = testData5[1399];
@(posedge clk);
#1;data_in = testData5[1400];
@(posedge clk);
#1;data_in = testData5[1401];
@(posedge clk);
#1;data_in = testData5[1402];
@(posedge clk);
#1;data_in = testData5[1403];
@(posedge clk);
#1;data_in = testData5[1404];
@(posedge clk);
#1;data_in = testData5[1405];
@(posedge clk);
#1;data_in = testData5[1406];
@(posedge clk);
#1;data_in = testData5[1407];
@(posedge clk);
#1;data_in = testData5[1408];
@(posedge clk);
#1;data_in = testData5[1409];
@(posedge clk);
#1;data_in = testData5[1410];
@(posedge clk);
#1;data_in = testData5[1411];
@(posedge clk);
#1;data_in = testData5[1412];
@(posedge clk);
#1;data_in = testData5[1413];
@(posedge clk);
#1;data_in = testData5[1414];
@(posedge clk);
#1;data_in = testData5[1415];
@(posedge clk);
#1;data_in = testData5[1416];
@(posedge clk);
#1;data_in = testData5[1417];
@(posedge clk);
#1;data_in = testData5[1418];
@(posedge clk);
#1;data_in = testData5[1419];
@(posedge clk);
#1;data_in = testData5[1420];
@(posedge clk);
#1;data_in = testData5[1421];
@(posedge clk);
#1;data_in = testData5[1422];
@(posedge clk);
#1;data_in = testData5[1423];
@(posedge clk);
#1;data_in = testData5[1424];
@(posedge clk);
#1;data_in = testData5[1425];
@(posedge clk);
#1;data_in = testData5[1426];
@(posedge clk);
#1;data_in = testData5[1427];
@(posedge clk);
#1;data_in = testData5[1428];
@(posedge clk);
#1;data_in = testData5[1429];
@(posedge clk);
#1;data_in = testData5[1430];
@(posedge clk);
#1;data_in = testData5[1431];
@(posedge clk);
#1;data_in = testData5[1432];
@(posedge clk);
#1;data_in = testData5[1433];
@(posedge clk);
#1;data_in = testData5[1434];
@(posedge clk);
#1;data_in = testData5[1435];
@(posedge clk);
#1;data_in = testData5[1436];
@(posedge clk);
#1;data_in = testData5[1437];
@(posedge clk);
#1;data_in = testData5[1438];
@(posedge clk);
#1;data_in = testData5[1439];
@(posedge clk);
#1;data_in = testData5[1440];
@(posedge clk);
#1;data_in = testData5[1441];
@(posedge clk);
#1;data_in = testData5[1442];
@(posedge clk);
#1;data_in = testData5[1443];
@(posedge clk);
#1;data_in = testData5[1444];
@(posedge clk);
#1;data_in = testData5[1445];
@(posedge clk);
#1;data_in = testData5[1446];
@(posedge clk);
#1;data_in = testData5[1447];
@(posedge clk);
#1;data_in = testData5[1448];
@(posedge clk);
#1;data_in = testData5[1449];
@(posedge clk);
#1;data_in = testData5[1450];
@(posedge clk);
#1;data_in = testData5[1451];
@(posedge clk);
#1;data_in = testData5[1452];
@(posedge clk);
#1;data_in = testData5[1453];
@(posedge clk);
#1;data_in = testData5[1454];
@(posedge clk);
#1;data_in = testData5[1455];
@(posedge clk);
#1;data_in = testData5[1456];
@(posedge clk);
#1;data_in = testData5[1457];
@(posedge clk);
#1;data_in = testData5[1458];
@(posedge clk);
#1;data_in = testData5[1459];
@(posedge clk);
#1;data_in = testData5[1460];
@(posedge clk);
#1;data_in = testData5[1461];
@(posedge clk);
#1;data_in = testData5[1462];
@(posedge clk);
#1;data_in = testData5[1463];
@(posedge clk);
#1;data_in = testData5[1464];
@(posedge clk);
#1;data_in = testData5[1465];
@(posedge clk);
#1;data_in = testData5[1466];
@(posedge clk);
#1;data_in = testData5[1467];
@(posedge clk);
#1;data_in = testData5[1468];
@(posedge clk);
#1;data_in = testData5[1469];
@(posedge clk);
#1;data_in = testData5[1470];
@(posedge clk);
#1;data_in = testData5[1471];
@(posedge clk);
#1;data_in = testData5[1472];
@(posedge clk);
#1;data_in = testData5[1473];
@(posedge clk);
#1;data_in = testData5[1474];
@(posedge clk);
#1;data_in = testData5[1475];
@(posedge clk);
#1;data_in = testData5[1476];
@(posedge clk);
#1;data_in = testData5[1477];
@(posedge clk);
#1;data_in = testData5[1478];
@(posedge clk);
#1;data_in = testData5[1479];
@(posedge clk);
#1;data_in = testData5[1480];
@(posedge clk);
#1;data_in = testData5[1481];
@(posedge clk);
#1;data_in = testData5[1482];
@(posedge clk);
#1;data_in = testData5[1483];
@(posedge clk);
#1;data_in = testData5[1484];
@(posedge clk);
#1;data_in = testData5[1485];
@(posedge clk);
#1;data_in = testData5[1486];
@(posedge clk);
#1;data_in = testData5[1487];
@(posedge clk);
#1;data_in = testData5[1488];
@(posedge clk);
#1;data_in = testData5[1489];
@(posedge clk);
#1;data_in = testData5[1490];
@(posedge clk);
#1;data_in = testData5[1491];
@(posedge clk);
#1;data_in = testData5[1492];
@(posedge clk);
#1;data_in = testData5[1493];
@(posedge clk);
#1;data_in = testData5[1494];
@(posedge clk);
#1;data_in = testData5[1495];
@(posedge clk);
#1;data_in = testData5[1496];
@(posedge clk);
#1;data_in = testData5[1497];
@(posedge clk);
#1;data_in = testData5[1498];
@(posedge clk);
#1;data_in = testData5[1499];
@(posedge clk);
#1;data_in = testData5[1500];
@(posedge clk);
#1;data_in = testData5[1501];
@(posedge clk);
#1;data_in = testData5[1502];
@(posedge clk);
#1;data_in = testData5[1503];
@(posedge clk);
#1;data_in = testData5[1504];
@(posedge clk);
#1;data_in = testData5[1505];
@(posedge clk);
#1;data_in = testData5[1506];
@(posedge clk);
#1;data_in = testData5[1507];
@(posedge clk);
#1;data_in = testData5[1508];
@(posedge clk);
#1;data_in = testData5[1509];
@(posedge clk);
#1;data_in = testData5[1510];
@(posedge clk);
#1;data_in = testData5[1511];
@(posedge clk);
#1;data_in = testData5[1512];
@(posedge clk);
#1;data_in = testData5[1513];
@(posedge clk);
#1;data_in = testData5[1514];
@(posedge clk);
#1;data_in = testData5[1515];
@(posedge clk);
#1;data_in = testData5[1516];
@(posedge clk);
#1;data_in = testData5[1517];
@(posedge clk);
#1;data_in = testData5[1518];
@(posedge clk);
#1;data_in = testData5[1519];
@(posedge clk);
#1;data_in = testData5[1520];
@(posedge clk);
#1;data_in = testData5[1521];
@(posedge clk);
#1;data_in = testData5[1522];
@(posedge clk);
#1;data_in = testData5[1523];
@(posedge clk);
#1;data_in = testData5[1524];
@(posedge clk);
#1;data_in = testData5[1525];
@(posedge clk);
#1;data_in = testData5[1526];
@(posedge clk);
#1;data_in = testData5[1527];
@(posedge clk);
#1;data_in = testData5[1528];
@(posedge clk);
#1;data_in = testData5[1529];
@(posedge clk);
#1;data_in = testData5[1530];
@(posedge clk);
#1;data_in = testData5[1531];
@(posedge clk);
#1;data_in = testData5[1532];
@(posedge clk);
#1;data_in = testData5[1533];
@(posedge clk);
#1;data_in = testData5[1534];
@(posedge clk);
#1;data_in = testData5[1535];
@(posedge clk);
#1;data_in = testData5[1536];
@(posedge clk);
#1;data_in = testData5[1537];
@(posedge clk);
#1;data_in = testData5[1538];
@(posedge clk);
#1;data_in = testData5[1539];
@(posedge clk);
#1;data_in = testData5[1540];
@(posedge clk);
#1;data_in = testData5[1541];
@(posedge clk);
#1;data_in = testData5[1542];
@(posedge clk);
#1;data_in = testData5[1543];
@(posedge clk);
#1;data_in = testData5[1544];
@(posedge clk);
#1;data_in = testData5[1545];
@(posedge clk);
#1;data_in = testData5[1546];
@(posedge clk);
#1;data_in = testData5[1547];
@(posedge clk);
#1;data_in = testData5[1548];
@(posedge clk);
#1;data_in = testData5[1549];
@(posedge clk);
#1;data_in = testData5[1550];
@(posedge clk);
#1;data_in = testData5[1551];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1552]; 
@(posedge clk);
#1;data_in = testData5[1553];
@(posedge clk);
#1;data_in = testData5[1554];
@(posedge clk);
#1;data_in = testData5[1555];
@(posedge clk);
#1;data_in = testData5[1556];
@(posedge clk);
#1;data_in = testData5[1557];
@(posedge clk);
#1;data_in = testData5[1558];
@(posedge clk);
#1;data_in = testData5[1559];
@(posedge clk);
#1;data_in = testData5[1560];
@(posedge clk);
#1;data_in = testData5[1561];
@(posedge clk);
#1;data_in = testData5[1562];
@(posedge clk);
#1;data_in = testData5[1563];
@(posedge clk);
#1;data_in = testData5[1564];
@(posedge clk);
#1;data_in = testData5[1565];
@(posedge clk);
#1;data_in = testData5[1566];
@(posedge clk);
#1;data_in = testData5[1567];
@(posedge clk);
#1;data_in = testData5[1568];
@(posedge clk);
#1;data_in = testData5[1569];
@(posedge clk);
#1;data_in = testData5[1570];
@(posedge clk);
#1;data_in = testData5[1571];
@(posedge clk);
#1;data_in = testData5[1572];
@(posedge clk);
#1;data_in = testData5[1573];
@(posedge clk);
#1;data_in = testData5[1574];
@(posedge clk);
#1;data_in = testData5[1575];
@(posedge clk);
#1;data_in = testData5[1576];
@(posedge clk);
#1;data_in = testData5[1577];
@(posedge clk);
#1;data_in = testData5[1578];
@(posedge clk);
#1;data_in = testData5[1579];
@(posedge clk);
#1;data_in = testData5[1580];
@(posedge clk);
#1;data_in = testData5[1581];
@(posedge clk);
#1;data_in = testData5[1582];
@(posedge clk);
#1;data_in = testData5[1583];
@(posedge clk);
#1;data_in = testData5[1584];
@(posedge clk);
#1;data_in = testData5[1585];
@(posedge clk);
#1;data_in = testData5[1586];
@(posedge clk);
#1;data_in = testData5[1587];
@(posedge clk);
#1;data_in = testData5[1588];
@(posedge clk);
#1;data_in = testData5[1589];
@(posedge clk);
#1;data_in = testData5[1590];
@(posedge clk);
#1;data_in = testData5[1591];
@(posedge clk);
#1;data_in = testData5[1592];
@(posedge clk);
#1;data_in = testData5[1593];
@(posedge clk);
#1;data_in = testData5[1594];
@(posedge clk);
#1;data_in = testData5[1595];
@(posedge clk);
#1;data_in = testData5[1596];
@(posedge clk);
#1;data_in = testData5[1597];
@(posedge clk);
#1;data_in = testData5[1598];
@(posedge clk);
#1;data_in = testData5[1599];
@(posedge clk);
#1;data_in = testData5[1600];
@(posedge clk);
#1;data_in = testData5[1601];
@(posedge clk);
#1;data_in = testData5[1602];
@(posedge clk);
#1;data_in = testData5[1603];
@(posedge clk);
#1;data_in = testData5[1604];
@(posedge clk);
#1;data_in = testData5[1605];
@(posedge clk);
#1;data_in = testData5[1606];
@(posedge clk);
#1;data_in = testData5[1607];
@(posedge clk);
#1;data_in = testData5[1608];
@(posedge clk);
#1;data_in = testData5[1609];
@(posedge clk);
#1;data_in = testData5[1610];
@(posedge clk);
#1;data_in = testData5[1611];
@(posedge clk);
#1;data_in = testData5[1612];
@(posedge clk);
#1;data_in = testData5[1613];
@(posedge clk);
#1;data_in = testData5[1614];
@(posedge clk);
#1;data_in = testData5[1615];
@(posedge clk);
#1;data_in = testData5[1616];
@(posedge clk);
#1;data_in = testData5[1617];
@(posedge clk);
#1;data_in = testData5[1618];
@(posedge clk);
#1;data_in = testData5[1619];
@(posedge clk);
#1;data_in = testData5[1620];
@(posedge clk);
#1;data_in = testData5[1621];
@(posedge clk);
#1;data_in = testData5[1622];
@(posedge clk);
#1;data_in = testData5[1623];
@(posedge clk);
#1;data_in = testData5[1624];
@(posedge clk);
#1;data_in = testData5[1625];
@(posedge clk);
#1;data_in = testData5[1626];
@(posedge clk);
#1;data_in = testData5[1627];
@(posedge clk);
#1;data_in = testData5[1628];
@(posedge clk);
#1;data_in = testData5[1629];
@(posedge clk);
#1;data_in = testData5[1630];
@(posedge clk);
#1;data_in = testData5[1631];
@(posedge clk);
#1;data_in = testData5[1632];
@(posedge clk);
#1;data_in = testData5[1633];
@(posedge clk);
#1;data_in = testData5[1634];
@(posedge clk);
#1;data_in = testData5[1635];
@(posedge clk);
#1;data_in = testData5[1636];
@(posedge clk);
#1;data_in = testData5[1637];
@(posedge clk);
#1;data_in = testData5[1638];
@(posedge clk);
#1;data_in = testData5[1639];
@(posedge clk);
#1;data_in = testData5[1640];
@(posedge clk);
#1;data_in = testData5[1641];
@(posedge clk);
#1;data_in = testData5[1642];
@(posedge clk);
#1;data_in = testData5[1643];
@(posedge clk);
#1;data_in = testData5[1644];
@(posedge clk);
#1;data_in = testData5[1645];
@(posedge clk);
#1;data_in = testData5[1646];
@(posedge clk);
#1;data_in = testData5[1647];
@(posedge clk);
#1;data_in = testData5[1648];
@(posedge clk);
#1;data_in = testData5[1649];
@(posedge clk);
#1;data_in = testData5[1650];
@(posedge clk);
#1;data_in = testData5[1651];
@(posedge clk);
#1;data_in = testData5[1652];
@(posedge clk);
#1;data_in = testData5[1653];
@(posedge clk);
#1;data_in = testData5[1654];
@(posedge clk);
#1;data_in = testData5[1655];
@(posedge clk);
#1;data_in = testData5[1656];
@(posedge clk);
#1;data_in = testData5[1657];
@(posedge clk);
#1;data_in = testData5[1658];
@(posedge clk);
#1;data_in = testData5[1659];
@(posedge clk);
#1;data_in = testData5[1660];
@(posedge clk);
#1;data_in = testData5[1661];
@(posedge clk);
#1;data_in = testData5[1662];
@(posedge clk);
#1;data_in = testData5[1663];
@(posedge clk);
#1;data_in = testData5[1664];
@(posedge clk);
#1;data_in = testData5[1665];
@(posedge clk);
#1;data_in = testData5[1666];
@(posedge clk);
#1;data_in = testData5[1667];
@(posedge clk);
#1;data_in = testData5[1668];
@(posedge clk);
#1;data_in = testData5[1669];
@(posedge clk);
#1;data_in = testData5[1670];
@(posedge clk);
#1;data_in = testData5[1671];
@(posedge clk);
#1;data_in = testData5[1672];
@(posedge clk);
#1;data_in = testData5[1673];
@(posedge clk);
#1;data_in = testData5[1674];
@(posedge clk);
#1;data_in = testData5[1675];
@(posedge clk);
#1;data_in = testData5[1676];
@(posedge clk);
#1;data_in = testData5[1677];
@(posedge clk);
#1;data_in = testData5[1678];
@(posedge clk);
#1;data_in = testData5[1679];
@(posedge clk);
#1;data_in = testData5[1680];
@(posedge clk);
#1;data_in = testData5[1681];
@(posedge clk);
#1;data_in = testData5[1682];
@(posedge clk);
#1;data_in = testData5[1683];
@(posedge clk);
#1;data_in = testData5[1684];
@(posedge clk);
#1;data_in = testData5[1685];
@(posedge clk);
#1;data_in = testData5[1686];
@(posedge clk);
#1;data_in = testData5[1687];
@(posedge clk);
#1;data_in = testData5[1688];
@(posedge clk);
#1;data_in = testData5[1689];
@(posedge clk);
#1;data_in = testData5[1690];
@(posedge clk);
#1;data_in = testData5[1691];
@(posedge clk);
#1;data_in = testData5[1692];
@(posedge clk);
#1;data_in = testData5[1693];
@(posedge clk);
#1;data_in = testData5[1694];
@(posedge clk);
#1;data_in = testData5[1695];
@(posedge clk);
#1;data_in = testData5[1696];
@(posedge clk);
#1;data_in = testData5[1697];
@(posedge clk);
#1;data_in = testData5[1698];
@(posedge clk);
#1;data_in = testData5[1699];
@(posedge clk);
#1;data_in = testData5[1700];
@(posedge clk);
#1;data_in = testData5[1701];
@(posedge clk);
#1;data_in = testData5[1702];
@(posedge clk);
#1;data_in = testData5[1703];
@(posedge clk);
#1;data_in = testData5[1704];
@(posedge clk);
#1;data_in = testData5[1705];
@(posedge clk);
#1;data_in = testData5[1706];
@(posedge clk);
#1;data_in = testData5[1707];
@(posedge clk);
#1;data_in = testData5[1708];
@(posedge clk);
#1;data_in = testData5[1709];
@(posedge clk);
#1;data_in = testData5[1710];
@(posedge clk);
#1;data_in = testData5[1711];
@(posedge clk);
#1;data_in = testData5[1712];
@(posedge clk);
#1;data_in = testData5[1713];
@(posedge clk);
#1;data_in = testData5[1714];
@(posedge clk);
#1;data_in = testData5[1715];
@(posedge clk);
#1;data_in = testData5[1716];
@(posedge clk);
#1;data_in = testData5[1717];
@(posedge clk);
#1;data_in = testData5[1718];
@(posedge clk);
#1;data_in = testData5[1719];
@(posedge clk);
#1;data_in = testData5[1720];
@(posedge clk);
#1;data_in = testData5[1721];
@(posedge clk);
#1;data_in = testData5[1722];
@(posedge clk);
#1;data_in = testData5[1723];
@(posedge clk);
#1;data_in = testData5[1724];
@(posedge clk);
#1;data_in = testData5[1725];
@(posedge clk);
#1;data_in = testData5[1726];
@(posedge clk);
#1;data_in = testData5[1727];
@(posedge clk);
#1;data_in = testData5[1728];
@(posedge clk);
#1;data_in = testData5[1729];
@(posedge clk);
#1;data_in = testData5[1730];
@(posedge clk);
#1;data_in = testData5[1731];
@(posedge clk);
#1;data_in = testData5[1732];
@(posedge clk);
#1;data_in = testData5[1733];
@(posedge clk);
#1;data_in = testData5[1734];
@(posedge clk);
#1;data_in = testData5[1735];
@(posedge clk);
#1;data_in = testData5[1736];
@(posedge clk);
#1;data_in = testData5[1737];
@(posedge clk);
#1;data_in = testData5[1738];
@(posedge clk);
#1;data_in = testData5[1739];
@(posedge clk);
#1;data_in = testData5[1740];
@(posedge clk);
#1;data_in = testData5[1741];
@(posedge clk);
#1;data_in = testData5[1742];
@(posedge clk);
#1;data_in = testData5[1743];
@(posedge clk);
#1;data_in = testData5[1744];
@(posedge clk);
#1;data_in = testData5[1745];
@(posedge clk);
#1;data_in = testData5[1746];
@(posedge clk);
#1;data_in = testData5[1747];
@(posedge clk);
#1;data_in = testData5[1748];
@(posedge clk);
#1;data_in = testData5[1749];
@(posedge clk);
#1;data_in = testData5[1750];
@(posedge clk);
#1;data_in = testData5[1751];
@(posedge clk);
#1;data_in = testData5[1752];
@(posedge clk);
#1;data_in = testData5[1753];
@(posedge clk);
#1;data_in = testData5[1754];
@(posedge clk);
#1;data_in = testData5[1755];
@(posedge clk);
#1;data_in = testData5[1756];
@(posedge clk);
#1;data_in = testData5[1757];
@(posedge clk);
#1;data_in = testData5[1758];
@(posedge clk);
#1;data_in = testData5[1759];
@(posedge clk);
#1;data_in = testData5[1760];
@(posedge clk);
#1;data_in = testData5[1761];
@(posedge clk);
#1;data_in = testData5[1762];
@(posedge clk);
#1;data_in = testData5[1763];
@(posedge clk);
#1;data_in = testData5[1764];
@(posedge clk);
#1;data_in = testData5[1765];
@(posedge clk);
#1;data_in = testData5[1766];
@(posedge clk);
#1;data_in = testData5[1767];
@(posedge clk);
#1;data_in = testData5[1768];
@(posedge clk);
#1;data_in = testData5[1769];
@(posedge clk);
#1;data_in = testData5[1770];
@(posedge clk);
#1;data_in = testData5[1771];
@(posedge clk);
#1;data_in = testData5[1772];
@(posedge clk);
#1;data_in = testData5[1773];
@(posedge clk);
#1;data_in = testData5[1774];
@(posedge clk);
#1;data_in = testData5[1775];
@(posedge clk);
#1;data_in = testData5[1776];
@(posedge clk);
#1;data_in = testData5[1777];
@(posedge clk);
#1;data_in = testData5[1778];
@(posedge clk);
#1;data_in = testData5[1779];
@(posedge clk);
#1;data_in = testData5[1780];
@(posedge clk);
#1;data_in = testData5[1781];
@(posedge clk);
#1;data_in = testData5[1782];
@(posedge clk);
#1;data_in = testData5[1783];
@(posedge clk);
#1;data_in = testData5[1784];
@(posedge clk);
#1;data_in = testData5[1785];
@(posedge clk);
#1;data_in = testData5[1786];
@(posedge clk);
#1;data_in = testData5[1787];
@(posedge clk);
#1;data_in = testData5[1788];
@(posedge clk);
#1;data_in = testData5[1789];
@(posedge clk);
#1;data_in = testData5[1790];
@(posedge clk);
#1;data_in = testData5[1791];
@(posedge clk);
#1;data_in = testData5[1792];
@(posedge clk);
#1;data_in = testData5[1793];
@(posedge clk);
#1;data_in = testData5[1794];
@(posedge clk);
#1;data_in = testData5[1795];
@(posedge clk);
#1;data_in = testData5[1796];
@(posedge clk);
#1;data_in = testData5[1797];
@(posedge clk);
#1;data_in = testData5[1798];
@(posedge clk);
#1;data_in = testData5[1799];
@(posedge clk);
#1;data_in = testData5[1800];
@(posedge clk);
#1;data_in = testData5[1801];
@(posedge clk);
#1;data_in = testData5[1802];
@(posedge clk);
#1;data_in = testData5[1803];
@(posedge clk);
#1;data_in = testData5[1804];
@(posedge clk);
#1;data_in = testData5[1805];
@(posedge clk);
#1;data_in = testData5[1806];
@(posedge clk);
#1;data_in = testData5[1807];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1808]; 
@(posedge clk);
#1;data_in = testData5[1809];
@(posedge clk);
#1;data_in = testData5[1810];
@(posedge clk);
#1;data_in = testData5[1811];
@(posedge clk);
#1;data_in = testData5[1812];
@(posedge clk);
#1;data_in = testData5[1813];
@(posedge clk);
#1;data_in = testData5[1814];
@(posedge clk);
#1;data_in = testData5[1815];
@(posedge clk);
#1;data_in = testData5[1816];
@(posedge clk);
#1;data_in = testData5[1817];
@(posedge clk);
#1;data_in = testData5[1818];
@(posedge clk);
#1;data_in = testData5[1819];
@(posedge clk);
#1;data_in = testData5[1820];
@(posedge clk);
#1;data_in = testData5[1821];
@(posedge clk);
#1;data_in = testData5[1822];
@(posedge clk);
#1;data_in = testData5[1823];
@(posedge clk);
#1;data_in = testData5[1824];
@(posedge clk);
#1;data_in = testData5[1825];
@(posedge clk);
#1;data_in = testData5[1826];
@(posedge clk);
#1;data_in = testData5[1827];
@(posedge clk);
#1;data_in = testData5[1828];
@(posedge clk);
#1;data_in = testData5[1829];
@(posedge clk);
#1;data_in = testData5[1830];
@(posedge clk);
#1;data_in = testData5[1831];
@(posedge clk);
#1;data_in = testData5[1832];
@(posedge clk);
#1;data_in = testData5[1833];
@(posedge clk);
#1;data_in = testData5[1834];
@(posedge clk);
#1;data_in = testData5[1835];
@(posedge clk);
#1;data_in = testData5[1836];
@(posedge clk);
#1;data_in = testData5[1837];
@(posedge clk);
#1;data_in = testData5[1838];
@(posedge clk);
#1;data_in = testData5[1839];
@(posedge clk);
#1;data_in = testData5[1840];
@(posedge clk);
#1;data_in = testData5[1841];
@(posedge clk);
#1;data_in = testData5[1842];
@(posedge clk);
#1;data_in = testData5[1843];
@(posedge clk);
#1;data_in = testData5[1844];
@(posedge clk);
#1;data_in = testData5[1845];
@(posedge clk);
#1;data_in = testData5[1846];
@(posedge clk);
#1;data_in = testData5[1847];
@(posedge clk);
#1;data_in = testData5[1848];
@(posedge clk);
#1;data_in = testData5[1849];
@(posedge clk);
#1;data_in = testData5[1850];
@(posedge clk);
#1;data_in = testData5[1851];
@(posedge clk);
#1;data_in = testData5[1852];
@(posedge clk);
#1;data_in = testData5[1853];
@(posedge clk);
#1;data_in = testData5[1854];
@(posedge clk);
#1;data_in = testData5[1855];
@(posedge clk);
#1;data_in = testData5[1856];
@(posedge clk);
#1;data_in = testData5[1857];
@(posedge clk);
#1;data_in = testData5[1858];
@(posedge clk);
#1;data_in = testData5[1859];
@(posedge clk);
#1;data_in = testData5[1860];
@(posedge clk);
#1;data_in = testData5[1861];
@(posedge clk);
#1;data_in = testData5[1862];
@(posedge clk);
#1;data_in = testData5[1863];
@(posedge clk);
#1;data_in = testData5[1864];
@(posedge clk);
#1;data_in = testData5[1865];
@(posedge clk);
#1;data_in = testData5[1866];
@(posedge clk);
#1;data_in = testData5[1867];
@(posedge clk);
#1;data_in = testData5[1868];
@(posedge clk);
#1;data_in = testData5[1869];
@(posedge clk);
#1;data_in = testData5[1870];
@(posedge clk);
#1;data_in = testData5[1871];
@(posedge clk);
#1;data_in = testData5[1872];
@(posedge clk);
#1;data_in = testData5[1873];
@(posedge clk);
#1;data_in = testData5[1874];
@(posedge clk);
#1;data_in = testData5[1875];
@(posedge clk);
#1;data_in = testData5[1876];
@(posedge clk);
#1;data_in = testData5[1877];
@(posedge clk);
#1;data_in = testData5[1878];
@(posedge clk);
#1;data_in = testData5[1879];
@(posedge clk);
#1;data_in = testData5[1880];
@(posedge clk);
#1;data_in = testData5[1881];
@(posedge clk);
#1;data_in = testData5[1882];
@(posedge clk);
#1;data_in = testData5[1883];
@(posedge clk);
#1;data_in = testData5[1884];
@(posedge clk);
#1;data_in = testData5[1885];
@(posedge clk);
#1;data_in = testData5[1886];
@(posedge clk);
#1;data_in = testData5[1887];
@(posedge clk);
#1;data_in = testData5[1888];
@(posedge clk);
#1;data_in = testData5[1889];
@(posedge clk);
#1;data_in = testData5[1890];
@(posedge clk);
#1;data_in = testData5[1891];
@(posedge clk);
#1;data_in = testData5[1892];
@(posedge clk);
#1;data_in = testData5[1893];
@(posedge clk);
#1;data_in = testData5[1894];
@(posedge clk);
#1;data_in = testData5[1895];
@(posedge clk);
#1;data_in = testData5[1896];
@(posedge clk);
#1;data_in = testData5[1897];
@(posedge clk);
#1;data_in = testData5[1898];
@(posedge clk);
#1;data_in = testData5[1899];
@(posedge clk);
#1;data_in = testData5[1900];
@(posedge clk);
#1;data_in = testData5[1901];
@(posedge clk);
#1;data_in = testData5[1902];
@(posedge clk);
#1;data_in = testData5[1903];
@(posedge clk);
#1;data_in = testData5[1904];
@(posedge clk);
#1;data_in = testData5[1905];
@(posedge clk);
#1;data_in = testData5[1906];
@(posedge clk);
#1;data_in = testData5[1907];
@(posedge clk);
#1;data_in = testData5[1908];
@(posedge clk);
#1;data_in = testData5[1909];
@(posedge clk);
#1;data_in = testData5[1910];
@(posedge clk);
#1;data_in = testData5[1911];
@(posedge clk);
#1;data_in = testData5[1912];
@(posedge clk);
#1;data_in = testData5[1913];
@(posedge clk);
#1;data_in = testData5[1914];
@(posedge clk);
#1;data_in = testData5[1915];
@(posedge clk);
#1;data_in = testData5[1916];
@(posedge clk);
#1;data_in = testData5[1917];
@(posedge clk);
#1;data_in = testData5[1918];
@(posedge clk);
#1;data_in = testData5[1919];
@(posedge clk);
#1;data_in = testData5[1920];
@(posedge clk);
#1;data_in = testData5[1921];
@(posedge clk);
#1;data_in = testData5[1922];
@(posedge clk);
#1;data_in = testData5[1923];
@(posedge clk);
#1;data_in = testData5[1924];
@(posedge clk);
#1;data_in = testData5[1925];
@(posedge clk);
#1;data_in = testData5[1926];
@(posedge clk);
#1;data_in = testData5[1927];
@(posedge clk);
#1;data_in = testData5[1928];
@(posedge clk);
#1;data_in = testData5[1929];
@(posedge clk);
#1;data_in = testData5[1930];
@(posedge clk);
#1;data_in = testData5[1931];
@(posedge clk);
#1;data_in = testData5[1932];
@(posedge clk);
#1;data_in = testData5[1933];
@(posedge clk);
#1;data_in = testData5[1934];
@(posedge clk);
#1;data_in = testData5[1935];
@(posedge clk);
#1;data_in = testData5[1936];
@(posedge clk);
#1;data_in = testData5[1937];
@(posedge clk);
#1;data_in = testData5[1938];
@(posedge clk);
#1;data_in = testData5[1939];
@(posedge clk);
#1;data_in = testData5[1940];
@(posedge clk);
#1;data_in = testData5[1941];
@(posedge clk);
#1;data_in = testData5[1942];
@(posedge clk);
#1;data_in = testData5[1943];
@(posedge clk);
#1;data_in = testData5[1944];
@(posedge clk);
#1;data_in = testData5[1945];
@(posedge clk);
#1;data_in = testData5[1946];
@(posedge clk);
#1;data_in = testData5[1947];
@(posedge clk);
#1;data_in = testData5[1948];
@(posedge clk);
#1;data_in = testData5[1949];
@(posedge clk);
#1;data_in = testData5[1950];
@(posedge clk);
#1;data_in = testData5[1951];
@(posedge clk);
#1;data_in = testData5[1952];
@(posedge clk);
#1;data_in = testData5[1953];
@(posedge clk);
#1;data_in = testData5[1954];
@(posedge clk);
#1;data_in = testData5[1955];
@(posedge clk);
#1;data_in = testData5[1956];
@(posedge clk);
#1;data_in = testData5[1957];
@(posedge clk);
#1;data_in = testData5[1958];
@(posedge clk);
#1;data_in = testData5[1959];
@(posedge clk);
#1;data_in = testData5[1960];
@(posedge clk);
#1;data_in = testData5[1961];
@(posedge clk);
#1;data_in = testData5[1962];
@(posedge clk);
#1;data_in = testData5[1963];
@(posedge clk);
#1;data_in = testData5[1964];
@(posedge clk);
#1;data_in = testData5[1965];
@(posedge clk);
#1;data_in = testData5[1966];
@(posedge clk);
#1;data_in = testData5[1967];
@(posedge clk);
#1;data_in = testData5[1968];
@(posedge clk);
#1;data_in = testData5[1969];
@(posedge clk);
#1;data_in = testData5[1970];
@(posedge clk);
#1;data_in = testData5[1971];
@(posedge clk);
#1;data_in = testData5[1972];
@(posedge clk);
#1;data_in = testData5[1973];
@(posedge clk);
#1;data_in = testData5[1974];
@(posedge clk);
#1;data_in = testData5[1975];
@(posedge clk);
#1;data_in = testData5[1976];
@(posedge clk);
#1;data_in = testData5[1977];
@(posedge clk);
#1;data_in = testData5[1978];
@(posedge clk);
#1;data_in = testData5[1979];
@(posedge clk);
#1;data_in = testData5[1980];
@(posedge clk);
#1;data_in = testData5[1981];
@(posedge clk);
#1;data_in = testData5[1982];
@(posedge clk);
#1;data_in = testData5[1983];
@(posedge clk);
#1;data_in = testData5[1984];
@(posedge clk);
#1;data_in = testData5[1985];
@(posedge clk);
#1;data_in = testData5[1986];
@(posedge clk);
#1;data_in = testData5[1987];
@(posedge clk);
#1;data_in = testData5[1988];
@(posedge clk);
#1;data_in = testData5[1989];
@(posedge clk);
#1;data_in = testData5[1990];
@(posedge clk);
#1;data_in = testData5[1991];
@(posedge clk);
#1;data_in = testData5[1992];
@(posedge clk);
#1;data_in = testData5[1993];
@(posedge clk);
#1;data_in = testData5[1994];
@(posedge clk);
#1;data_in = testData5[1995];
@(posedge clk);
#1;data_in = testData5[1996];
@(posedge clk);
#1;data_in = testData5[1997];
@(posedge clk);
#1;data_in = testData5[1998];
@(posedge clk);
#1;data_in = testData5[1999];
@(posedge clk);
#1;data_in = testData5[2000];
@(posedge clk);
#1;data_in = testData5[2001];
@(posedge clk);
#1;data_in = testData5[2002];
@(posedge clk);
#1;data_in = testData5[2003];
@(posedge clk);
#1;data_in = testData5[2004];
@(posedge clk);
#1;data_in = testData5[2005];
@(posedge clk);
#1;data_in = testData5[2006];
@(posedge clk);
#1;data_in = testData5[2007];
@(posedge clk);
#1;data_in = testData5[2008];
@(posedge clk);
#1;data_in = testData5[2009];
@(posedge clk);
#1;data_in = testData5[2010];
@(posedge clk);
#1;data_in = testData5[2011];
@(posedge clk);
#1;data_in = testData5[2012];
@(posedge clk);
#1;data_in = testData5[2013];
@(posedge clk);
#1;data_in = testData5[2014];
@(posedge clk);
#1;data_in = testData5[2015];
@(posedge clk);
#1;data_in = testData5[2016];
@(posedge clk);
#1;data_in = testData5[2017];
@(posedge clk);
#1;data_in = testData5[2018];
@(posedge clk);
#1;data_in = testData5[2019];
@(posedge clk);
#1;data_in = testData5[2020];
@(posedge clk);
#1;data_in = testData5[2021];
@(posedge clk);
#1;data_in = testData5[2022];
@(posedge clk);
#1;data_in = testData5[2023];
@(posedge clk);
#1;data_in = testData5[2024];
@(posedge clk);
#1;data_in = testData5[2025];
@(posedge clk);
#1;data_in = testData5[2026];
@(posedge clk);
#1;data_in = testData5[2027];
@(posedge clk);
#1;data_in = testData5[2028];
@(posedge clk);
#1;data_in = testData5[2029];
@(posedge clk);
#1;data_in = testData5[2030];
@(posedge clk);
#1;data_in = testData5[2031];
@(posedge clk);
#1;data_in = testData5[2032];
@(posedge clk);
#1;data_in = testData5[2033];
@(posedge clk);
#1;data_in = testData5[2034];
@(posedge clk);
#1;data_in = testData5[2035];
@(posedge clk);
#1;data_in = testData5[2036];
@(posedge clk);
#1;data_in = testData5[2037];
@(posedge clk);
#1;data_in = testData5[2038];
@(posedge clk);
#1;data_in = testData5[2039];
@(posedge clk);
#1;data_in = testData5[2040];
@(posedge clk);
#1;data_in = testData5[2041];
@(posedge clk);
#1;data_in = testData5[2042];
@(posedge clk);
#1;data_in = testData5[2043];
@(posedge clk);
#1;data_in = testData5[2044];
@(posedge clk);
#1;data_in = testData5[2045];
@(posedge clk);
#1;data_in = testData5[2046];
@(posedge clk);
#1;data_in = testData5[2047];
@(posedge clk);
#1;data_in = testData5[2048];
@(posedge clk);
#1;data_in = testData5[2049];
@(posedge clk);
#1;data_in = testData5[2050];
@(posedge clk);
#1;data_in = testData5[2051];
@(posedge clk);
#1;data_in = testData5[2052];
@(posedge clk);
#1;data_in = testData5[2053];
@(posedge clk);
#1;data_in = testData5[2054];
@(posedge clk);
#1;data_in = testData5[2055];
@(posedge clk);
#1;data_in = testData5[2056];
@(posedge clk);
#1;data_in = testData5[2057];
@(posedge clk);
#1;data_in = testData5[2058];
@(posedge clk);
#1;data_in = testData5[2059];
@(posedge clk);
#1;data_in = testData5[2060];
@(posedge clk);
#1;data_in = testData5[2061];
@(posedge clk);
#1;data_in = testData5[2062];
@(posedge clk);
#1;data_in = testData5[2063];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2064]; 
@(posedge clk);
#1;data_in = testData5[2065];
@(posedge clk);
#1;data_in = testData5[2066];
@(posedge clk);
#1;data_in = testData5[2067];
@(posedge clk);
#1;data_in = testData5[2068];
@(posedge clk);
#1;data_in = testData5[2069];
@(posedge clk);
#1;data_in = testData5[2070];
@(posedge clk);
#1;data_in = testData5[2071];
@(posedge clk);
#1;data_in = testData5[2072];
@(posedge clk);
#1;data_in = testData5[2073];
@(posedge clk);
#1;data_in = testData5[2074];
@(posedge clk);
#1;data_in = testData5[2075];
@(posedge clk);
#1;data_in = testData5[2076];
@(posedge clk);
#1;data_in = testData5[2077];
@(posedge clk);
#1;data_in = testData5[2078];
@(posedge clk);
#1;data_in = testData5[2079];
@(posedge clk);
#1;data_in = testData5[2080];
@(posedge clk);
#1;data_in = testData5[2081];
@(posedge clk);
#1;data_in = testData5[2082];
@(posedge clk);
#1;data_in = testData5[2083];
@(posedge clk);
#1;data_in = testData5[2084];
@(posedge clk);
#1;data_in = testData5[2085];
@(posedge clk);
#1;data_in = testData5[2086];
@(posedge clk);
#1;data_in = testData5[2087];
@(posedge clk);
#1;data_in = testData5[2088];
@(posedge clk);
#1;data_in = testData5[2089];
@(posedge clk);
#1;data_in = testData5[2090];
@(posedge clk);
#1;data_in = testData5[2091];
@(posedge clk);
#1;data_in = testData5[2092];
@(posedge clk);
#1;data_in = testData5[2093];
@(posedge clk);
#1;data_in = testData5[2094];
@(posedge clk);
#1;data_in = testData5[2095];
@(posedge clk);
#1;data_in = testData5[2096];
@(posedge clk);
#1;data_in = testData5[2097];
@(posedge clk);
#1;data_in = testData5[2098];
@(posedge clk);
#1;data_in = testData5[2099];
@(posedge clk);
#1;data_in = testData5[2100];
@(posedge clk);
#1;data_in = testData5[2101];
@(posedge clk);
#1;data_in = testData5[2102];
@(posedge clk);
#1;data_in = testData5[2103];
@(posedge clk);
#1;data_in = testData5[2104];
@(posedge clk);
#1;data_in = testData5[2105];
@(posedge clk);
#1;data_in = testData5[2106];
@(posedge clk);
#1;data_in = testData5[2107];
@(posedge clk);
#1;data_in = testData5[2108];
@(posedge clk);
#1;data_in = testData5[2109];
@(posedge clk);
#1;data_in = testData5[2110];
@(posedge clk);
#1;data_in = testData5[2111];
@(posedge clk);
#1;data_in = testData5[2112];
@(posedge clk);
#1;data_in = testData5[2113];
@(posedge clk);
#1;data_in = testData5[2114];
@(posedge clk);
#1;data_in = testData5[2115];
@(posedge clk);
#1;data_in = testData5[2116];
@(posedge clk);
#1;data_in = testData5[2117];
@(posedge clk);
#1;data_in = testData5[2118];
@(posedge clk);
#1;data_in = testData5[2119];
@(posedge clk);
#1;data_in = testData5[2120];
@(posedge clk);
#1;data_in = testData5[2121];
@(posedge clk);
#1;data_in = testData5[2122];
@(posedge clk);
#1;data_in = testData5[2123];
@(posedge clk);
#1;data_in = testData5[2124];
@(posedge clk);
#1;data_in = testData5[2125];
@(posedge clk);
#1;data_in = testData5[2126];
@(posedge clk);
#1;data_in = testData5[2127];
@(posedge clk);
#1;data_in = testData5[2128];
@(posedge clk);
#1;data_in = testData5[2129];
@(posedge clk);
#1;data_in = testData5[2130];
@(posedge clk);
#1;data_in = testData5[2131];
@(posedge clk);
#1;data_in = testData5[2132];
@(posedge clk);
#1;data_in = testData5[2133];
@(posedge clk);
#1;data_in = testData5[2134];
@(posedge clk);
#1;data_in = testData5[2135];
@(posedge clk);
#1;data_in = testData5[2136];
@(posedge clk);
#1;data_in = testData5[2137];
@(posedge clk);
#1;data_in = testData5[2138];
@(posedge clk);
#1;data_in = testData5[2139];
@(posedge clk);
#1;data_in = testData5[2140];
@(posedge clk);
#1;data_in = testData5[2141];
@(posedge clk);
#1;data_in = testData5[2142];
@(posedge clk);
#1;data_in = testData5[2143];
@(posedge clk);
#1;data_in = testData5[2144];
@(posedge clk);
#1;data_in = testData5[2145];
@(posedge clk);
#1;data_in = testData5[2146];
@(posedge clk);
#1;data_in = testData5[2147];
@(posedge clk);
#1;data_in = testData5[2148];
@(posedge clk);
#1;data_in = testData5[2149];
@(posedge clk);
#1;data_in = testData5[2150];
@(posedge clk);
#1;data_in = testData5[2151];
@(posedge clk);
#1;data_in = testData5[2152];
@(posedge clk);
#1;data_in = testData5[2153];
@(posedge clk);
#1;data_in = testData5[2154];
@(posedge clk);
#1;data_in = testData5[2155];
@(posedge clk);
#1;data_in = testData5[2156];
@(posedge clk);
#1;data_in = testData5[2157];
@(posedge clk);
#1;data_in = testData5[2158];
@(posedge clk);
#1;data_in = testData5[2159];
@(posedge clk);
#1;data_in = testData5[2160];
@(posedge clk);
#1;data_in = testData5[2161];
@(posedge clk);
#1;data_in = testData5[2162];
@(posedge clk);
#1;data_in = testData5[2163];
@(posedge clk);
#1;data_in = testData5[2164];
@(posedge clk);
#1;data_in = testData5[2165];
@(posedge clk);
#1;data_in = testData5[2166];
@(posedge clk);
#1;data_in = testData5[2167];
@(posedge clk);
#1;data_in = testData5[2168];
@(posedge clk);
#1;data_in = testData5[2169];
@(posedge clk);
#1;data_in = testData5[2170];
@(posedge clk);
#1;data_in = testData5[2171];
@(posedge clk);
#1;data_in = testData5[2172];
@(posedge clk);
#1;data_in = testData5[2173];
@(posedge clk);
#1;data_in = testData5[2174];
@(posedge clk);
#1;data_in = testData5[2175];
@(posedge clk);
#1;data_in = testData5[2176];
@(posedge clk);
#1;data_in = testData5[2177];
@(posedge clk);
#1;data_in = testData5[2178];
@(posedge clk);
#1;data_in = testData5[2179];
@(posedge clk);
#1;data_in = testData5[2180];
@(posedge clk);
#1;data_in = testData5[2181];
@(posedge clk);
#1;data_in = testData5[2182];
@(posedge clk);
#1;data_in = testData5[2183];
@(posedge clk);
#1;data_in = testData5[2184];
@(posedge clk);
#1;data_in = testData5[2185];
@(posedge clk);
#1;data_in = testData5[2186];
@(posedge clk);
#1;data_in = testData5[2187];
@(posedge clk);
#1;data_in = testData5[2188];
@(posedge clk);
#1;data_in = testData5[2189];
@(posedge clk);
#1;data_in = testData5[2190];
@(posedge clk);
#1;data_in = testData5[2191];
@(posedge clk);
#1;data_in = testData5[2192];
@(posedge clk);
#1;data_in = testData5[2193];
@(posedge clk);
#1;data_in = testData5[2194];
@(posedge clk);
#1;data_in = testData5[2195];
@(posedge clk);
#1;data_in = testData5[2196];
@(posedge clk);
#1;data_in = testData5[2197];
@(posedge clk);
#1;data_in = testData5[2198];
@(posedge clk);
#1;data_in = testData5[2199];
@(posedge clk);
#1;data_in = testData5[2200];
@(posedge clk);
#1;data_in = testData5[2201];
@(posedge clk);
#1;data_in = testData5[2202];
@(posedge clk);
#1;data_in = testData5[2203];
@(posedge clk);
#1;data_in = testData5[2204];
@(posedge clk);
#1;data_in = testData5[2205];
@(posedge clk);
#1;data_in = testData5[2206];
@(posedge clk);
#1;data_in = testData5[2207];
@(posedge clk);
#1;data_in = testData5[2208];
@(posedge clk);
#1;data_in = testData5[2209];
@(posedge clk);
#1;data_in = testData5[2210];
@(posedge clk);
#1;data_in = testData5[2211];
@(posedge clk);
#1;data_in = testData5[2212];
@(posedge clk);
#1;data_in = testData5[2213];
@(posedge clk);
#1;data_in = testData5[2214];
@(posedge clk);
#1;data_in = testData5[2215];
@(posedge clk);
#1;data_in = testData5[2216];
@(posedge clk);
#1;data_in = testData5[2217];
@(posedge clk);
#1;data_in = testData5[2218];
@(posedge clk);
#1;data_in = testData5[2219];
@(posedge clk);
#1;data_in = testData5[2220];
@(posedge clk);
#1;data_in = testData5[2221];
@(posedge clk);
#1;data_in = testData5[2222];
@(posedge clk);
#1;data_in = testData5[2223];
@(posedge clk);
#1;data_in = testData5[2224];
@(posedge clk);
#1;data_in = testData5[2225];
@(posedge clk);
#1;data_in = testData5[2226];
@(posedge clk);
#1;data_in = testData5[2227];
@(posedge clk);
#1;data_in = testData5[2228];
@(posedge clk);
#1;data_in = testData5[2229];
@(posedge clk);
#1;data_in = testData5[2230];
@(posedge clk);
#1;data_in = testData5[2231];
@(posedge clk);
#1;data_in = testData5[2232];
@(posedge clk);
#1;data_in = testData5[2233];
@(posedge clk);
#1;data_in = testData5[2234];
@(posedge clk);
#1;data_in = testData5[2235];
@(posedge clk);
#1;data_in = testData5[2236];
@(posedge clk);
#1;data_in = testData5[2237];
@(posedge clk);
#1;data_in = testData5[2238];
@(posedge clk);
#1;data_in = testData5[2239];
@(posedge clk);
#1;data_in = testData5[2240];
@(posedge clk);
#1;data_in = testData5[2241];
@(posedge clk);
#1;data_in = testData5[2242];
@(posedge clk);
#1;data_in = testData5[2243];
@(posedge clk);
#1;data_in = testData5[2244];
@(posedge clk);
#1;data_in = testData5[2245];
@(posedge clk);
#1;data_in = testData5[2246];
@(posedge clk);
#1;data_in = testData5[2247];
@(posedge clk);
#1;data_in = testData5[2248];
@(posedge clk);
#1;data_in = testData5[2249];
@(posedge clk);
#1;data_in = testData5[2250];
@(posedge clk);
#1;data_in = testData5[2251];
@(posedge clk);
#1;data_in = testData5[2252];
@(posedge clk);
#1;data_in = testData5[2253];
@(posedge clk);
#1;data_in = testData5[2254];
@(posedge clk);
#1;data_in = testData5[2255];
@(posedge clk);
#1;data_in = testData5[2256];
@(posedge clk);
#1;data_in = testData5[2257];
@(posedge clk);
#1;data_in = testData5[2258];
@(posedge clk);
#1;data_in = testData5[2259];
@(posedge clk);
#1;data_in = testData5[2260];
@(posedge clk);
#1;data_in = testData5[2261];
@(posedge clk);
#1;data_in = testData5[2262];
@(posedge clk);
#1;data_in = testData5[2263];
@(posedge clk);
#1;data_in = testData5[2264];
@(posedge clk);
#1;data_in = testData5[2265];
@(posedge clk);
#1;data_in = testData5[2266];
@(posedge clk);
#1;data_in = testData5[2267];
@(posedge clk);
#1;data_in = testData5[2268];
@(posedge clk);
#1;data_in = testData5[2269];
@(posedge clk);
#1;data_in = testData5[2270];
@(posedge clk);
#1;data_in = testData5[2271];
@(posedge clk);
#1;data_in = testData5[2272];
@(posedge clk);
#1;data_in = testData5[2273];
@(posedge clk);
#1;data_in = testData5[2274];
@(posedge clk);
#1;data_in = testData5[2275];
@(posedge clk);
#1;data_in = testData5[2276];
@(posedge clk);
#1;data_in = testData5[2277];
@(posedge clk);
#1;data_in = testData5[2278];
@(posedge clk);
#1;data_in = testData5[2279];
@(posedge clk);
#1;data_in = testData5[2280];
@(posedge clk);
#1;data_in = testData5[2281];
@(posedge clk);
#1;data_in = testData5[2282];
@(posedge clk);
#1;data_in = testData5[2283];
@(posedge clk);
#1;data_in = testData5[2284];
@(posedge clk);
#1;data_in = testData5[2285];
@(posedge clk);
#1;data_in = testData5[2286];
@(posedge clk);
#1;data_in = testData5[2287];
@(posedge clk);
#1;data_in = testData5[2288];
@(posedge clk);
#1;data_in = testData5[2289];
@(posedge clk);
#1;data_in = testData5[2290];
@(posedge clk);
#1;data_in = testData5[2291];
@(posedge clk);
#1;data_in = testData5[2292];
@(posedge clk);
#1;data_in = testData5[2293];
@(posedge clk);
#1;data_in = testData5[2294];
@(posedge clk);
#1;data_in = testData5[2295];
@(posedge clk);
#1;data_in = testData5[2296];
@(posedge clk);
#1;data_in = testData5[2297];
@(posedge clk);
#1;data_in = testData5[2298];
@(posedge clk);
#1;data_in = testData5[2299];
@(posedge clk);
#1;data_in = testData5[2300];
@(posedge clk);
#1;data_in = testData5[2301];
@(posedge clk);
#1;data_in = testData5[2302];
@(posedge clk);
#1;data_in = testData5[2303];
@(posedge clk);
#1;data_in = testData5[2304];
@(posedge clk);
#1;data_in = testData5[2305];
@(posedge clk);
#1;data_in = testData5[2306];
@(posedge clk);
#1;data_in = testData5[2307];
@(posedge clk);
#1;data_in = testData5[2308];
@(posedge clk);
#1;data_in = testData5[2309];
@(posedge clk);
#1;data_in = testData5[2310];
@(posedge clk);
#1;data_in = testData5[2311];
@(posedge clk);
#1;data_in = testData5[2312];
@(posedge clk);
#1;data_in = testData5[2313];
@(posedge clk);
#1;data_in = testData5[2314];
@(posedge clk);
#1;data_in = testData5[2315];
@(posedge clk);
#1;data_in = testData5[2316];
@(posedge clk);
#1;data_in = testData5[2317];
@(posedge clk);
#1;data_in = testData5[2318];
@(posedge clk);
#1;data_in = testData5[2319];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2320]; 
@(posedge clk);
#1;data_in = testData5[2321];
@(posedge clk);
#1;data_in = testData5[2322];
@(posedge clk);
#1;data_in = testData5[2323];
@(posedge clk);
#1;data_in = testData5[2324];
@(posedge clk);
#1;data_in = testData5[2325];
@(posedge clk);
#1;data_in = testData5[2326];
@(posedge clk);
#1;data_in = testData5[2327];
@(posedge clk);
#1;data_in = testData5[2328];
@(posedge clk);
#1;data_in = testData5[2329];
@(posedge clk);
#1;data_in = testData5[2330];
@(posedge clk);
#1;data_in = testData5[2331];
@(posedge clk);
#1;data_in = testData5[2332];
@(posedge clk);
#1;data_in = testData5[2333];
@(posedge clk);
#1;data_in = testData5[2334];
@(posedge clk);
#1;data_in = testData5[2335];
@(posedge clk);
#1;data_in = testData5[2336];
@(posedge clk);
#1;data_in = testData5[2337];
@(posedge clk);
#1;data_in = testData5[2338];
@(posedge clk);
#1;data_in = testData5[2339];
@(posedge clk);
#1;data_in = testData5[2340];
@(posedge clk);
#1;data_in = testData5[2341];
@(posedge clk);
#1;data_in = testData5[2342];
@(posedge clk);
#1;data_in = testData5[2343];
@(posedge clk);
#1;data_in = testData5[2344];
@(posedge clk);
#1;data_in = testData5[2345];
@(posedge clk);
#1;data_in = testData5[2346];
@(posedge clk);
#1;data_in = testData5[2347];
@(posedge clk);
#1;data_in = testData5[2348];
@(posedge clk);
#1;data_in = testData5[2349];
@(posedge clk);
#1;data_in = testData5[2350];
@(posedge clk);
#1;data_in = testData5[2351];
@(posedge clk);
#1;data_in = testData5[2352];
@(posedge clk);
#1;data_in = testData5[2353];
@(posedge clk);
#1;data_in = testData5[2354];
@(posedge clk);
#1;data_in = testData5[2355];
@(posedge clk);
#1;data_in = testData5[2356];
@(posedge clk);
#1;data_in = testData5[2357];
@(posedge clk);
#1;data_in = testData5[2358];
@(posedge clk);
#1;data_in = testData5[2359];
@(posedge clk);
#1;data_in = testData5[2360];
@(posedge clk);
#1;data_in = testData5[2361];
@(posedge clk);
#1;data_in = testData5[2362];
@(posedge clk);
#1;data_in = testData5[2363];
@(posedge clk);
#1;data_in = testData5[2364];
@(posedge clk);
#1;data_in = testData5[2365];
@(posedge clk);
#1;data_in = testData5[2366];
@(posedge clk);
#1;data_in = testData5[2367];
@(posedge clk);
#1;data_in = testData5[2368];
@(posedge clk);
#1;data_in = testData5[2369];
@(posedge clk);
#1;data_in = testData5[2370];
@(posedge clk);
#1;data_in = testData5[2371];
@(posedge clk);
#1;data_in = testData5[2372];
@(posedge clk);
#1;data_in = testData5[2373];
@(posedge clk);
#1;data_in = testData5[2374];
@(posedge clk);
#1;data_in = testData5[2375];
@(posedge clk);
#1;data_in = testData5[2376];
@(posedge clk);
#1;data_in = testData5[2377];
@(posedge clk);
#1;data_in = testData5[2378];
@(posedge clk);
#1;data_in = testData5[2379];
@(posedge clk);
#1;data_in = testData5[2380];
@(posedge clk);
#1;data_in = testData5[2381];
@(posedge clk);
#1;data_in = testData5[2382];
@(posedge clk);
#1;data_in = testData5[2383];
@(posedge clk);
#1;data_in = testData5[2384];
@(posedge clk);
#1;data_in = testData5[2385];
@(posedge clk);
#1;data_in = testData5[2386];
@(posedge clk);
#1;data_in = testData5[2387];
@(posedge clk);
#1;data_in = testData5[2388];
@(posedge clk);
#1;data_in = testData5[2389];
@(posedge clk);
#1;data_in = testData5[2390];
@(posedge clk);
#1;data_in = testData5[2391];
@(posedge clk);
#1;data_in = testData5[2392];
@(posedge clk);
#1;data_in = testData5[2393];
@(posedge clk);
#1;data_in = testData5[2394];
@(posedge clk);
#1;data_in = testData5[2395];
@(posedge clk);
#1;data_in = testData5[2396];
@(posedge clk);
#1;data_in = testData5[2397];
@(posedge clk);
#1;data_in = testData5[2398];
@(posedge clk);
#1;data_in = testData5[2399];
@(posedge clk);
#1;data_in = testData5[2400];
@(posedge clk);
#1;data_in = testData5[2401];
@(posedge clk);
#1;data_in = testData5[2402];
@(posedge clk);
#1;data_in = testData5[2403];
@(posedge clk);
#1;data_in = testData5[2404];
@(posedge clk);
#1;data_in = testData5[2405];
@(posedge clk);
#1;data_in = testData5[2406];
@(posedge clk);
#1;data_in = testData5[2407];
@(posedge clk);
#1;data_in = testData5[2408];
@(posedge clk);
#1;data_in = testData5[2409];
@(posedge clk);
#1;data_in = testData5[2410];
@(posedge clk);
#1;data_in = testData5[2411];
@(posedge clk);
#1;data_in = testData5[2412];
@(posedge clk);
#1;data_in = testData5[2413];
@(posedge clk);
#1;data_in = testData5[2414];
@(posedge clk);
#1;data_in = testData5[2415];
@(posedge clk);
#1;data_in = testData5[2416];
@(posedge clk);
#1;data_in = testData5[2417];
@(posedge clk);
#1;data_in = testData5[2418];
@(posedge clk);
#1;data_in = testData5[2419];
@(posedge clk);
#1;data_in = testData5[2420];
@(posedge clk);
#1;data_in = testData5[2421];
@(posedge clk);
#1;data_in = testData5[2422];
@(posedge clk);
#1;data_in = testData5[2423];
@(posedge clk);
#1;data_in = testData5[2424];
@(posedge clk);
#1;data_in = testData5[2425];
@(posedge clk);
#1;data_in = testData5[2426];
@(posedge clk);
#1;data_in = testData5[2427];
@(posedge clk);
#1;data_in = testData5[2428];
@(posedge clk);
#1;data_in = testData5[2429];
@(posedge clk);
#1;data_in = testData5[2430];
@(posedge clk);
#1;data_in = testData5[2431];
@(posedge clk);
#1;data_in = testData5[2432];
@(posedge clk);
#1;data_in = testData5[2433];
@(posedge clk);
#1;data_in = testData5[2434];
@(posedge clk);
#1;data_in = testData5[2435];
@(posedge clk);
#1;data_in = testData5[2436];
@(posedge clk);
#1;data_in = testData5[2437];
@(posedge clk);
#1;data_in = testData5[2438];
@(posedge clk);
#1;data_in = testData5[2439];
@(posedge clk);
#1;data_in = testData5[2440];
@(posedge clk);
#1;data_in = testData5[2441];
@(posedge clk);
#1;data_in = testData5[2442];
@(posedge clk);
#1;data_in = testData5[2443];
@(posedge clk);
#1;data_in = testData5[2444];
@(posedge clk);
#1;data_in = testData5[2445];
@(posedge clk);
#1;data_in = testData5[2446];
@(posedge clk);
#1;data_in = testData5[2447];
@(posedge clk);
#1;data_in = testData5[2448];
@(posedge clk);
#1;data_in = testData5[2449];
@(posedge clk);
#1;data_in = testData5[2450];
@(posedge clk);
#1;data_in = testData5[2451];
@(posedge clk);
#1;data_in = testData5[2452];
@(posedge clk);
#1;data_in = testData5[2453];
@(posedge clk);
#1;data_in = testData5[2454];
@(posedge clk);
#1;data_in = testData5[2455];
@(posedge clk);
#1;data_in = testData5[2456];
@(posedge clk);
#1;data_in = testData5[2457];
@(posedge clk);
#1;data_in = testData5[2458];
@(posedge clk);
#1;data_in = testData5[2459];
@(posedge clk);
#1;data_in = testData5[2460];
@(posedge clk);
#1;data_in = testData5[2461];
@(posedge clk);
#1;data_in = testData5[2462];
@(posedge clk);
#1;data_in = testData5[2463];
@(posedge clk);
#1;data_in = testData5[2464];
@(posedge clk);
#1;data_in = testData5[2465];
@(posedge clk);
#1;data_in = testData5[2466];
@(posedge clk);
#1;data_in = testData5[2467];
@(posedge clk);
#1;data_in = testData5[2468];
@(posedge clk);
#1;data_in = testData5[2469];
@(posedge clk);
#1;data_in = testData5[2470];
@(posedge clk);
#1;data_in = testData5[2471];
@(posedge clk);
#1;data_in = testData5[2472];
@(posedge clk);
#1;data_in = testData5[2473];
@(posedge clk);
#1;data_in = testData5[2474];
@(posedge clk);
#1;data_in = testData5[2475];
@(posedge clk);
#1;data_in = testData5[2476];
@(posedge clk);
#1;data_in = testData5[2477];
@(posedge clk);
#1;data_in = testData5[2478];
@(posedge clk);
#1;data_in = testData5[2479];
@(posedge clk);
#1;data_in = testData5[2480];
@(posedge clk);
#1;data_in = testData5[2481];
@(posedge clk);
#1;data_in = testData5[2482];
@(posedge clk);
#1;data_in = testData5[2483];
@(posedge clk);
#1;data_in = testData5[2484];
@(posedge clk);
#1;data_in = testData5[2485];
@(posedge clk);
#1;data_in = testData5[2486];
@(posedge clk);
#1;data_in = testData5[2487];
@(posedge clk);
#1;data_in = testData5[2488];
@(posedge clk);
#1;data_in = testData5[2489];
@(posedge clk);
#1;data_in = testData5[2490];
@(posedge clk);
#1;data_in = testData5[2491];
@(posedge clk);
#1;data_in = testData5[2492];
@(posedge clk);
#1;data_in = testData5[2493];
@(posedge clk);
#1;data_in = testData5[2494];
@(posedge clk);
#1;data_in = testData5[2495];
@(posedge clk);
#1;data_in = testData5[2496];
@(posedge clk);
#1;data_in = testData5[2497];
@(posedge clk);
#1;data_in = testData5[2498];
@(posedge clk);
#1;data_in = testData5[2499];
@(posedge clk);
#1;data_in = testData5[2500];
@(posedge clk);
#1;data_in = testData5[2501];
@(posedge clk);
#1;data_in = testData5[2502];
@(posedge clk);
#1;data_in = testData5[2503];
@(posedge clk);
#1;data_in = testData5[2504];
@(posedge clk);
#1;data_in = testData5[2505];
@(posedge clk);
#1;data_in = testData5[2506];
@(posedge clk);
#1;data_in = testData5[2507];
@(posedge clk);
#1;data_in = testData5[2508];
@(posedge clk);
#1;data_in = testData5[2509];
@(posedge clk);
#1;data_in = testData5[2510];
@(posedge clk);
#1;data_in = testData5[2511];
@(posedge clk);
#1;data_in = testData5[2512];
@(posedge clk);
#1;data_in = testData5[2513];
@(posedge clk);
#1;data_in = testData5[2514];
@(posedge clk);
#1;data_in = testData5[2515];
@(posedge clk);
#1;data_in = testData5[2516];
@(posedge clk);
#1;data_in = testData5[2517];
@(posedge clk);
#1;data_in = testData5[2518];
@(posedge clk);
#1;data_in = testData5[2519];
@(posedge clk);
#1;data_in = testData5[2520];
@(posedge clk);
#1;data_in = testData5[2521];
@(posedge clk);
#1;data_in = testData5[2522];
@(posedge clk);
#1;data_in = testData5[2523];
@(posedge clk);
#1;data_in = testData5[2524];
@(posedge clk);
#1;data_in = testData5[2525];
@(posedge clk);
#1;data_in = testData5[2526];
@(posedge clk);
#1;data_in = testData5[2527];
@(posedge clk);
#1;data_in = testData5[2528];
@(posedge clk);
#1;data_in = testData5[2529];
@(posedge clk);
#1;data_in = testData5[2530];
@(posedge clk);
#1;data_in = testData5[2531];
@(posedge clk);
#1;data_in = testData5[2532];
@(posedge clk);
#1;data_in = testData5[2533];
@(posedge clk);
#1;data_in = testData5[2534];
@(posedge clk);
#1;data_in = testData5[2535];
@(posedge clk);
#1;data_in = testData5[2536];
@(posedge clk);
#1;data_in = testData5[2537];
@(posedge clk);
#1;data_in = testData5[2538];
@(posedge clk);
#1;data_in = testData5[2539];
@(posedge clk);
#1;data_in = testData5[2540];
@(posedge clk);
#1;data_in = testData5[2541];
@(posedge clk);
#1;data_in = testData5[2542];
@(posedge clk);
#1;data_in = testData5[2543];
@(posedge clk);
#1;data_in = testData5[2544];
@(posedge clk);
#1;data_in = testData5[2545];
@(posedge clk);
#1;data_in = testData5[2546];
@(posedge clk);
#1;data_in = testData5[2547];
@(posedge clk);
#1;data_in = testData5[2548];
@(posedge clk);
#1;data_in = testData5[2549];
@(posedge clk);
#1;data_in = testData5[2550];
@(posedge clk);
#1;data_in = testData5[2551];
@(posedge clk);
#1;data_in = testData5[2552];
@(posedge clk);
#1;data_in = testData5[2553];
@(posedge clk);
#1;data_in = testData5[2554];
@(posedge clk);
#1;data_in = testData5[2555];
@(posedge clk);
#1;data_in = testData5[2556];
@(posedge clk);
#1;data_in = testData5[2557];
@(posedge clk);
#1;data_in = testData5[2558];
@(posedge clk);
#1;data_in = testData5[2559];
@(posedge clk);
#1;data_in = testData5[2560];
@(posedge clk);
#1;data_in = testData5[2561];
@(posedge clk);
#1;data_in = testData5[2562];
@(posedge clk);
#1;data_in = testData5[2563];
@(posedge clk);
#1;data_in = testData5[2564];
@(posedge clk);
#1;data_in = testData5[2565];
@(posedge clk);
#1;data_in = testData5[2566];
@(posedge clk);
#1;data_in = testData5[2567];
@(posedge clk);
#1;data_in = testData5[2568];
@(posedge clk);
#1;data_in = testData5[2569];
@(posedge clk);
#1;data_in = testData5[2570];
@(posedge clk);
#1;data_in = testData5[2571];
@(posedge clk);
#1;data_in = testData5[2572];
@(posedge clk);
#1;data_in = testData5[2573];
@(posedge clk);
#1;data_in = testData5[2574];
@(posedge clk);
#1;data_in = testData5[2575];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2576]; 
@(posedge clk);
#1;data_in = testData5[2577];
@(posedge clk);
#1;data_in = testData5[2578];
@(posedge clk);
#1;data_in = testData5[2579];
@(posedge clk);
#1;data_in = testData5[2580];
@(posedge clk);
#1;data_in = testData5[2581];
@(posedge clk);
#1;data_in = testData5[2582];
@(posedge clk);
#1;data_in = testData5[2583];
@(posedge clk);
#1;data_in = testData5[2584];
@(posedge clk);
#1;data_in = testData5[2585];
@(posedge clk);
#1;data_in = testData5[2586];
@(posedge clk);
#1;data_in = testData5[2587];
@(posedge clk);
#1;data_in = testData5[2588];
@(posedge clk);
#1;data_in = testData5[2589];
@(posedge clk);
#1;data_in = testData5[2590];
@(posedge clk);
#1;data_in = testData5[2591];
@(posedge clk);
#1;data_in = testData5[2592];
@(posedge clk);
#1;data_in = testData5[2593];
@(posedge clk);
#1;data_in = testData5[2594];
@(posedge clk);
#1;data_in = testData5[2595];
@(posedge clk);
#1;data_in = testData5[2596];
@(posedge clk);
#1;data_in = testData5[2597];
@(posedge clk);
#1;data_in = testData5[2598];
@(posedge clk);
#1;data_in = testData5[2599];
@(posedge clk);
#1;data_in = testData5[2600];
@(posedge clk);
#1;data_in = testData5[2601];
@(posedge clk);
#1;data_in = testData5[2602];
@(posedge clk);
#1;data_in = testData5[2603];
@(posedge clk);
#1;data_in = testData5[2604];
@(posedge clk);
#1;data_in = testData5[2605];
@(posedge clk);
#1;data_in = testData5[2606];
@(posedge clk);
#1;data_in = testData5[2607];
@(posedge clk);
#1;data_in = testData5[2608];
@(posedge clk);
#1;data_in = testData5[2609];
@(posedge clk);
#1;data_in = testData5[2610];
@(posedge clk);
#1;data_in = testData5[2611];
@(posedge clk);
#1;data_in = testData5[2612];
@(posedge clk);
#1;data_in = testData5[2613];
@(posedge clk);
#1;data_in = testData5[2614];
@(posedge clk);
#1;data_in = testData5[2615];
@(posedge clk);
#1;data_in = testData5[2616];
@(posedge clk);
#1;data_in = testData5[2617];
@(posedge clk);
#1;data_in = testData5[2618];
@(posedge clk);
#1;data_in = testData5[2619];
@(posedge clk);
#1;data_in = testData5[2620];
@(posedge clk);
#1;data_in = testData5[2621];
@(posedge clk);
#1;data_in = testData5[2622];
@(posedge clk);
#1;data_in = testData5[2623];
@(posedge clk);
#1;data_in = testData5[2624];
@(posedge clk);
#1;data_in = testData5[2625];
@(posedge clk);
#1;data_in = testData5[2626];
@(posedge clk);
#1;data_in = testData5[2627];
@(posedge clk);
#1;data_in = testData5[2628];
@(posedge clk);
#1;data_in = testData5[2629];
@(posedge clk);
#1;data_in = testData5[2630];
@(posedge clk);
#1;data_in = testData5[2631];
@(posedge clk);
#1;data_in = testData5[2632];
@(posedge clk);
#1;data_in = testData5[2633];
@(posedge clk);
#1;data_in = testData5[2634];
@(posedge clk);
#1;data_in = testData5[2635];
@(posedge clk);
#1;data_in = testData5[2636];
@(posedge clk);
#1;data_in = testData5[2637];
@(posedge clk);
#1;data_in = testData5[2638];
@(posedge clk);
#1;data_in = testData5[2639];
@(posedge clk);
#1;data_in = testData5[2640];
@(posedge clk);
#1;data_in = testData5[2641];
@(posedge clk);
#1;data_in = testData5[2642];
@(posedge clk);
#1;data_in = testData5[2643];
@(posedge clk);
#1;data_in = testData5[2644];
@(posedge clk);
#1;data_in = testData5[2645];
@(posedge clk);
#1;data_in = testData5[2646];
@(posedge clk);
#1;data_in = testData5[2647];
@(posedge clk);
#1;data_in = testData5[2648];
@(posedge clk);
#1;data_in = testData5[2649];
@(posedge clk);
#1;data_in = testData5[2650];
@(posedge clk);
#1;data_in = testData5[2651];
@(posedge clk);
#1;data_in = testData5[2652];
@(posedge clk);
#1;data_in = testData5[2653];
@(posedge clk);
#1;data_in = testData5[2654];
@(posedge clk);
#1;data_in = testData5[2655];
@(posedge clk);
#1;data_in = testData5[2656];
@(posedge clk);
#1;data_in = testData5[2657];
@(posedge clk);
#1;data_in = testData5[2658];
@(posedge clk);
#1;data_in = testData5[2659];
@(posedge clk);
#1;data_in = testData5[2660];
@(posedge clk);
#1;data_in = testData5[2661];
@(posedge clk);
#1;data_in = testData5[2662];
@(posedge clk);
#1;data_in = testData5[2663];
@(posedge clk);
#1;data_in = testData5[2664];
@(posedge clk);
#1;data_in = testData5[2665];
@(posedge clk);
#1;data_in = testData5[2666];
@(posedge clk);
#1;data_in = testData5[2667];
@(posedge clk);
#1;data_in = testData5[2668];
@(posedge clk);
#1;data_in = testData5[2669];
@(posedge clk);
#1;data_in = testData5[2670];
@(posedge clk);
#1;data_in = testData5[2671];
@(posedge clk);
#1;data_in = testData5[2672];
@(posedge clk);
#1;data_in = testData5[2673];
@(posedge clk);
#1;data_in = testData5[2674];
@(posedge clk);
#1;data_in = testData5[2675];
@(posedge clk);
#1;data_in = testData5[2676];
@(posedge clk);
#1;data_in = testData5[2677];
@(posedge clk);
#1;data_in = testData5[2678];
@(posedge clk);
#1;data_in = testData5[2679];
@(posedge clk);
#1;data_in = testData5[2680];
@(posedge clk);
#1;data_in = testData5[2681];
@(posedge clk);
#1;data_in = testData5[2682];
@(posedge clk);
#1;data_in = testData5[2683];
@(posedge clk);
#1;data_in = testData5[2684];
@(posedge clk);
#1;data_in = testData5[2685];
@(posedge clk);
#1;data_in = testData5[2686];
@(posedge clk);
#1;data_in = testData5[2687];
@(posedge clk);
#1;data_in = testData5[2688];
@(posedge clk);
#1;data_in = testData5[2689];
@(posedge clk);
#1;data_in = testData5[2690];
@(posedge clk);
#1;data_in = testData5[2691];
@(posedge clk);
#1;data_in = testData5[2692];
@(posedge clk);
#1;data_in = testData5[2693];
@(posedge clk);
#1;data_in = testData5[2694];
@(posedge clk);
#1;data_in = testData5[2695];
@(posedge clk);
#1;data_in = testData5[2696];
@(posedge clk);
#1;data_in = testData5[2697];
@(posedge clk);
#1;data_in = testData5[2698];
@(posedge clk);
#1;data_in = testData5[2699];
@(posedge clk);
#1;data_in = testData5[2700];
@(posedge clk);
#1;data_in = testData5[2701];
@(posedge clk);
#1;data_in = testData5[2702];
@(posedge clk);
#1;data_in = testData5[2703];
@(posedge clk);
#1;data_in = testData5[2704];
@(posedge clk);
#1;data_in = testData5[2705];
@(posedge clk);
#1;data_in = testData5[2706];
@(posedge clk);
#1;data_in = testData5[2707];
@(posedge clk);
#1;data_in = testData5[2708];
@(posedge clk);
#1;data_in = testData5[2709];
@(posedge clk);
#1;data_in = testData5[2710];
@(posedge clk);
#1;data_in = testData5[2711];
@(posedge clk);
#1;data_in = testData5[2712];
@(posedge clk);
#1;data_in = testData5[2713];
@(posedge clk);
#1;data_in = testData5[2714];
@(posedge clk);
#1;data_in = testData5[2715];
@(posedge clk);
#1;data_in = testData5[2716];
@(posedge clk);
#1;data_in = testData5[2717];
@(posedge clk);
#1;data_in = testData5[2718];
@(posedge clk);
#1;data_in = testData5[2719];
@(posedge clk);
#1;data_in = testData5[2720];
@(posedge clk);
#1;data_in = testData5[2721];
@(posedge clk);
#1;data_in = testData5[2722];
@(posedge clk);
#1;data_in = testData5[2723];
@(posedge clk);
#1;data_in = testData5[2724];
@(posedge clk);
#1;data_in = testData5[2725];
@(posedge clk);
#1;data_in = testData5[2726];
@(posedge clk);
#1;data_in = testData5[2727];
@(posedge clk);
#1;data_in = testData5[2728];
@(posedge clk);
#1;data_in = testData5[2729];
@(posedge clk);
#1;data_in = testData5[2730];
@(posedge clk);
#1;data_in = testData5[2731];
@(posedge clk);
#1;data_in = testData5[2732];
@(posedge clk);
#1;data_in = testData5[2733];
@(posedge clk);
#1;data_in = testData5[2734];
@(posedge clk);
#1;data_in = testData5[2735];
@(posedge clk);
#1;data_in = testData5[2736];
@(posedge clk);
#1;data_in = testData5[2737];
@(posedge clk);
#1;data_in = testData5[2738];
@(posedge clk);
#1;data_in = testData5[2739];
@(posedge clk);
#1;data_in = testData5[2740];
@(posedge clk);
#1;data_in = testData5[2741];
@(posedge clk);
#1;data_in = testData5[2742];
@(posedge clk);
#1;data_in = testData5[2743];
@(posedge clk);
#1;data_in = testData5[2744];
@(posedge clk);
#1;data_in = testData5[2745];
@(posedge clk);
#1;data_in = testData5[2746];
@(posedge clk);
#1;data_in = testData5[2747];
@(posedge clk);
#1;data_in = testData5[2748];
@(posedge clk);
#1;data_in = testData5[2749];
@(posedge clk);
#1;data_in = testData5[2750];
@(posedge clk);
#1;data_in = testData5[2751];
@(posedge clk);
#1;data_in = testData5[2752];
@(posedge clk);
#1;data_in = testData5[2753];
@(posedge clk);
#1;data_in = testData5[2754];
@(posedge clk);
#1;data_in = testData5[2755];
@(posedge clk);
#1;data_in = testData5[2756];
@(posedge clk);
#1;data_in = testData5[2757];
@(posedge clk);
#1;data_in = testData5[2758];
@(posedge clk);
#1;data_in = testData5[2759];
@(posedge clk);
#1;data_in = testData5[2760];
@(posedge clk);
#1;data_in = testData5[2761];
@(posedge clk);
#1;data_in = testData5[2762];
@(posedge clk);
#1;data_in = testData5[2763];
@(posedge clk);
#1;data_in = testData5[2764];
@(posedge clk);
#1;data_in = testData5[2765];
@(posedge clk);
#1;data_in = testData5[2766];
@(posedge clk);
#1;data_in = testData5[2767];
@(posedge clk);
#1;data_in = testData5[2768];
@(posedge clk);
#1;data_in = testData5[2769];
@(posedge clk);
#1;data_in = testData5[2770];
@(posedge clk);
#1;data_in = testData5[2771];
@(posedge clk);
#1;data_in = testData5[2772];
@(posedge clk);
#1;data_in = testData5[2773];
@(posedge clk);
#1;data_in = testData5[2774];
@(posedge clk);
#1;data_in = testData5[2775];
@(posedge clk);
#1;data_in = testData5[2776];
@(posedge clk);
#1;data_in = testData5[2777];
@(posedge clk);
#1;data_in = testData5[2778];
@(posedge clk);
#1;data_in = testData5[2779];
@(posedge clk);
#1;data_in = testData5[2780];
@(posedge clk);
#1;data_in = testData5[2781];
@(posedge clk);
#1;data_in = testData5[2782];
@(posedge clk);
#1;data_in = testData5[2783];
@(posedge clk);
#1;data_in = testData5[2784];
@(posedge clk);
#1;data_in = testData5[2785];
@(posedge clk);
#1;data_in = testData5[2786];
@(posedge clk);
#1;data_in = testData5[2787];
@(posedge clk);
#1;data_in = testData5[2788];
@(posedge clk);
#1;data_in = testData5[2789];
@(posedge clk);
#1;data_in = testData5[2790];
@(posedge clk);
#1;data_in = testData5[2791];
@(posedge clk);
#1;data_in = testData5[2792];
@(posedge clk);
#1;data_in = testData5[2793];
@(posedge clk);
#1;data_in = testData5[2794];
@(posedge clk);
#1;data_in = testData5[2795];
@(posedge clk);
#1;data_in = testData5[2796];
@(posedge clk);
#1;data_in = testData5[2797];
@(posedge clk);
#1;data_in = testData5[2798];
@(posedge clk);
#1;data_in = testData5[2799];
@(posedge clk);
#1;data_in = testData5[2800];
@(posedge clk);
#1;data_in = testData5[2801];
@(posedge clk);
#1;data_in = testData5[2802];
@(posedge clk);
#1;data_in = testData5[2803];
@(posedge clk);
#1;data_in = testData5[2804];
@(posedge clk);
#1;data_in = testData5[2805];
@(posedge clk);
#1;data_in = testData5[2806];
@(posedge clk);
#1;data_in = testData5[2807];
@(posedge clk);
#1;data_in = testData5[2808];
@(posedge clk);
#1;data_in = testData5[2809];
@(posedge clk);
#1;data_in = testData5[2810];
@(posedge clk);
#1;data_in = testData5[2811];
@(posedge clk);
#1;data_in = testData5[2812];
@(posedge clk);
#1;data_in = testData5[2813];
@(posedge clk);
#1;data_in = testData5[2814];
@(posedge clk);
#1;data_in = testData5[2815];
@(posedge clk);
#1;data_in = testData5[2816];
@(posedge clk);
#1;data_in = testData5[2817];
@(posedge clk);
#1;data_in = testData5[2818];
@(posedge clk);
#1;data_in = testData5[2819];
@(posedge clk);
#1;data_in = testData5[2820];
@(posedge clk);
#1;data_in = testData5[2821];
@(posedge clk);
#1;data_in = testData5[2822];
@(posedge clk);
#1;data_in = testData5[2823];
@(posedge clk);
#1;data_in = testData5[2824];
@(posedge clk);
#1;data_in = testData5[2825];
@(posedge clk);
#1;data_in = testData5[2826];
@(posedge clk);
#1;data_in = testData5[2827];
@(posedge clk);
#1;data_in = testData5[2828];
@(posedge clk);
#1;data_in = testData5[2829];
@(posedge clk);
#1;data_in = testData5[2830];
@(posedge clk);
#1;data_in = testData5[2831];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2832]; 
@(posedge clk);
#1;data_in = testData5[2833];
@(posedge clk);
#1;data_in = testData5[2834];
@(posedge clk);
#1;data_in = testData5[2835];
@(posedge clk);
#1;data_in = testData5[2836];
@(posedge clk);
#1;data_in = testData5[2837];
@(posedge clk);
#1;data_in = testData5[2838];
@(posedge clk);
#1;data_in = testData5[2839];
@(posedge clk);
#1;data_in = testData5[2840];
@(posedge clk);
#1;data_in = testData5[2841];
@(posedge clk);
#1;data_in = testData5[2842];
@(posedge clk);
#1;data_in = testData5[2843];
@(posedge clk);
#1;data_in = testData5[2844];
@(posedge clk);
#1;data_in = testData5[2845];
@(posedge clk);
#1;data_in = testData5[2846];
@(posedge clk);
#1;data_in = testData5[2847];
@(posedge clk);
#1;data_in = testData5[2848];
@(posedge clk);
#1;data_in = testData5[2849];
@(posedge clk);
#1;data_in = testData5[2850];
@(posedge clk);
#1;data_in = testData5[2851];
@(posedge clk);
#1;data_in = testData5[2852];
@(posedge clk);
#1;data_in = testData5[2853];
@(posedge clk);
#1;data_in = testData5[2854];
@(posedge clk);
#1;data_in = testData5[2855];
@(posedge clk);
#1;data_in = testData5[2856];
@(posedge clk);
#1;data_in = testData5[2857];
@(posedge clk);
#1;data_in = testData5[2858];
@(posedge clk);
#1;data_in = testData5[2859];
@(posedge clk);
#1;data_in = testData5[2860];
@(posedge clk);
#1;data_in = testData5[2861];
@(posedge clk);
#1;data_in = testData5[2862];
@(posedge clk);
#1;data_in = testData5[2863];
@(posedge clk);
#1;data_in = testData5[2864];
@(posedge clk);
#1;data_in = testData5[2865];
@(posedge clk);
#1;data_in = testData5[2866];
@(posedge clk);
#1;data_in = testData5[2867];
@(posedge clk);
#1;data_in = testData5[2868];
@(posedge clk);
#1;data_in = testData5[2869];
@(posedge clk);
#1;data_in = testData5[2870];
@(posedge clk);
#1;data_in = testData5[2871];
@(posedge clk);
#1;data_in = testData5[2872];
@(posedge clk);
#1;data_in = testData5[2873];
@(posedge clk);
#1;data_in = testData5[2874];
@(posedge clk);
#1;data_in = testData5[2875];
@(posedge clk);
#1;data_in = testData5[2876];
@(posedge clk);
#1;data_in = testData5[2877];
@(posedge clk);
#1;data_in = testData5[2878];
@(posedge clk);
#1;data_in = testData5[2879];
@(posedge clk);
#1;data_in = testData5[2880];
@(posedge clk);
#1;data_in = testData5[2881];
@(posedge clk);
#1;data_in = testData5[2882];
@(posedge clk);
#1;data_in = testData5[2883];
@(posedge clk);
#1;data_in = testData5[2884];
@(posedge clk);
#1;data_in = testData5[2885];
@(posedge clk);
#1;data_in = testData5[2886];
@(posedge clk);
#1;data_in = testData5[2887];
@(posedge clk);
#1;data_in = testData5[2888];
@(posedge clk);
#1;data_in = testData5[2889];
@(posedge clk);
#1;data_in = testData5[2890];
@(posedge clk);
#1;data_in = testData5[2891];
@(posedge clk);
#1;data_in = testData5[2892];
@(posedge clk);
#1;data_in = testData5[2893];
@(posedge clk);
#1;data_in = testData5[2894];
@(posedge clk);
#1;data_in = testData5[2895];
@(posedge clk);
#1;data_in = testData5[2896];
@(posedge clk);
#1;data_in = testData5[2897];
@(posedge clk);
#1;data_in = testData5[2898];
@(posedge clk);
#1;data_in = testData5[2899];
@(posedge clk);
#1;data_in = testData5[2900];
@(posedge clk);
#1;data_in = testData5[2901];
@(posedge clk);
#1;data_in = testData5[2902];
@(posedge clk);
#1;data_in = testData5[2903];
@(posedge clk);
#1;data_in = testData5[2904];
@(posedge clk);
#1;data_in = testData5[2905];
@(posedge clk);
#1;data_in = testData5[2906];
@(posedge clk);
#1;data_in = testData5[2907];
@(posedge clk);
#1;data_in = testData5[2908];
@(posedge clk);
#1;data_in = testData5[2909];
@(posedge clk);
#1;data_in = testData5[2910];
@(posedge clk);
#1;data_in = testData5[2911];
@(posedge clk);
#1;data_in = testData5[2912];
@(posedge clk);
#1;data_in = testData5[2913];
@(posedge clk);
#1;data_in = testData5[2914];
@(posedge clk);
#1;data_in = testData5[2915];
@(posedge clk);
#1;data_in = testData5[2916];
@(posedge clk);
#1;data_in = testData5[2917];
@(posedge clk);
#1;data_in = testData5[2918];
@(posedge clk);
#1;data_in = testData5[2919];
@(posedge clk);
#1;data_in = testData5[2920];
@(posedge clk);
#1;data_in = testData5[2921];
@(posedge clk);
#1;data_in = testData5[2922];
@(posedge clk);
#1;data_in = testData5[2923];
@(posedge clk);
#1;data_in = testData5[2924];
@(posedge clk);
#1;data_in = testData5[2925];
@(posedge clk);
#1;data_in = testData5[2926];
@(posedge clk);
#1;data_in = testData5[2927];
@(posedge clk);
#1;data_in = testData5[2928];
@(posedge clk);
#1;data_in = testData5[2929];
@(posedge clk);
#1;data_in = testData5[2930];
@(posedge clk);
#1;data_in = testData5[2931];
@(posedge clk);
#1;data_in = testData5[2932];
@(posedge clk);
#1;data_in = testData5[2933];
@(posedge clk);
#1;data_in = testData5[2934];
@(posedge clk);
#1;data_in = testData5[2935];
@(posedge clk);
#1;data_in = testData5[2936];
@(posedge clk);
#1;data_in = testData5[2937];
@(posedge clk);
#1;data_in = testData5[2938];
@(posedge clk);
#1;data_in = testData5[2939];
@(posedge clk);
#1;data_in = testData5[2940];
@(posedge clk);
#1;data_in = testData5[2941];
@(posedge clk);
#1;data_in = testData5[2942];
@(posedge clk);
#1;data_in = testData5[2943];
@(posedge clk);
#1;data_in = testData5[2944];
@(posedge clk);
#1;data_in = testData5[2945];
@(posedge clk);
#1;data_in = testData5[2946];
@(posedge clk);
#1;data_in = testData5[2947];
@(posedge clk);
#1;data_in = testData5[2948];
@(posedge clk);
#1;data_in = testData5[2949];
@(posedge clk);
#1;data_in = testData5[2950];
@(posedge clk);
#1;data_in = testData5[2951];
@(posedge clk);
#1;data_in = testData5[2952];
@(posedge clk);
#1;data_in = testData5[2953];
@(posedge clk);
#1;data_in = testData5[2954];
@(posedge clk);
#1;data_in = testData5[2955];
@(posedge clk);
#1;data_in = testData5[2956];
@(posedge clk);
#1;data_in = testData5[2957];
@(posedge clk);
#1;data_in = testData5[2958];
@(posedge clk);
#1;data_in = testData5[2959];
@(posedge clk);
#1;data_in = testData5[2960];
@(posedge clk);
#1;data_in = testData5[2961];
@(posedge clk);
#1;data_in = testData5[2962];
@(posedge clk);
#1;data_in = testData5[2963];
@(posedge clk);
#1;data_in = testData5[2964];
@(posedge clk);
#1;data_in = testData5[2965];
@(posedge clk);
#1;data_in = testData5[2966];
@(posedge clk);
#1;data_in = testData5[2967];
@(posedge clk);
#1;data_in = testData5[2968];
@(posedge clk);
#1;data_in = testData5[2969];
@(posedge clk);
#1;data_in = testData5[2970];
@(posedge clk);
#1;data_in = testData5[2971];
@(posedge clk);
#1;data_in = testData5[2972];
@(posedge clk);
#1;data_in = testData5[2973];
@(posedge clk);
#1;data_in = testData5[2974];
@(posedge clk);
#1;data_in = testData5[2975];
@(posedge clk);
#1;data_in = testData5[2976];
@(posedge clk);
#1;data_in = testData5[2977];
@(posedge clk);
#1;data_in = testData5[2978];
@(posedge clk);
#1;data_in = testData5[2979];
@(posedge clk);
#1;data_in = testData5[2980];
@(posedge clk);
#1;data_in = testData5[2981];
@(posedge clk);
#1;data_in = testData5[2982];
@(posedge clk);
#1;data_in = testData5[2983];
@(posedge clk);
#1;data_in = testData5[2984];
@(posedge clk);
#1;data_in = testData5[2985];
@(posedge clk);
#1;data_in = testData5[2986];
@(posedge clk);
#1;data_in = testData5[2987];
@(posedge clk);
#1;data_in = testData5[2988];
@(posedge clk);
#1;data_in = testData5[2989];
@(posedge clk);
#1;data_in = testData5[2990];
@(posedge clk);
#1;data_in = testData5[2991];
@(posedge clk);
#1;data_in = testData5[2992];
@(posedge clk);
#1;data_in = testData5[2993];
@(posedge clk);
#1;data_in = testData5[2994];
@(posedge clk);
#1;data_in = testData5[2995];
@(posedge clk);
#1;data_in = testData5[2996];
@(posedge clk);
#1;data_in = testData5[2997];
@(posedge clk);
#1;data_in = testData5[2998];
@(posedge clk);
#1;data_in = testData5[2999];
@(posedge clk);
#1;data_in = testData5[3000];
@(posedge clk);
#1;data_in = testData5[3001];
@(posedge clk);
#1;data_in = testData5[3002];
@(posedge clk);
#1;data_in = testData5[3003];
@(posedge clk);
#1;data_in = testData5[3004];
@(posedge clk);
#1;data_in = testData5[3005];
@(posedge clk);
#1;data_in = testData5[3006];
@(posedge clk);
#1;data_in = testData5[3007];
@(posedge clk);
#1;data_in = testData5[3008];
@(posedge clk);
#1;data_in = testData5[3009];
@(posedge clk);
#1;data_in = testData5[3010];
@(posedge clk);
#1;data_in = testData5[3011];
@(posedge clk);
#1;data_in = testData5[3012];
@(posedge clk);
#1;data_in = testData5[3013];
@(posedge clk);
#1;data_in = testData5[3014];
@(posedge clk);
#1;data_in = testData5[3015];
@(posedge clk);
#1;data_in = testData5[3016];
@(posedge clk);
#1;data_in = testData5[3017];
@(posedge clk);
#1;data_in = testData5[3018];
@(posedge clk);
#1;data_in = testData5[3019];
@(posedge clk);
#1;data_in = testData5[3020];
@(posedge clk);
#1;data_in = testData5[3021];
@(posedge clk);
#1;data_in = testData5[3022];
@(posedge clk);
#1;data_in = testData5[3023];
@(posedge clk);
#1;data_in = testData5[3024];
@(posedge clk);
#1;data_in = testData5[3025];
@(posedge clk);
#1;data_in = testData5[3026];
@(posedge clk);
#1;data_in = testData5[3027];
@(posedge clk);
#1;data_in = testData5[3028];
@(posedge clk);
#1;data_in = testData5[3029];
@(posedge clk);
#1;data_in = testData5[3030];
@(posedge clk);
#1;data_in = testData5[3031];
@(posedge clk);
#1;data_in = testData5[3032];
@(posedge clk);
#1;data_in = testData5[3033];
@(posedge clk);
#1;data_in = testData5[3034];
@(posedge clk);
#1;data_in = testData5[3035];
@(posedge clk);
#1;data_in = testData5[3036];
@(posedge clk);
#1;data_in = testData5[3037];
@(posedge clk);
#1;data_in = testData5[3038];
@(posedge clk);
#1;data_in = testData5[3039];
@(posedge clk);
#1;data_in = testData5[3040];
@(posedge clk);
#1;data_in = testData5[3041];
@(posedge clk);
#1;data_in = testData5[3042];
@(posedge clk);
#1;data_in = testData5[3043];
@(posedge clk);
#1;data_in = testData5[3044];
@(posedge clk);
#1;data_in = testData5[3045];
@(posedge clk);
#1;data_in = testData5[3046];
@(posedge clk);
#1;data_in = testData5[3047];
@(posedge clk);
#1;data_in = testData5[3048];
@(posedge clk);
#1;data_in = testData5[3049];
@(posedge clk);
#1;data_in = testData5[3050];
@(posedge clk);
#1;data_in = testData5[3051];
@(posedge clk);
#1;data_in = testData5[3052];
@(posedge clk);
#1;data_in = testData5[3053];
@(posedge clk);
#1;data_in = testData5[3054];
@(posedge clk);
#1;data_in = testData5[3055];
@(posedge clk);
#1;data_in = testData5[3056];
@(posedge clk);
#1;data_in = testData5[3057];
@(posedge clk);
#1;data_in = testData5[3058];
@(posedge clk);
#1;data_in = testData5[3059];
@(posedge clk);
#1;data_in = testData5[3060];
@(posedge clk);
#1;data_in = testData5[3061];
@(posedge clk);
#1;data_in = testData5[3062];
@(posedge clk);
#1;data_in = testData5[3063];
@(posedge clk);
#1;data_in = testData5[3064];
@(posedge clk);
#1;data_in = testData5[3065];
@(posedge clk);
#1;data_in = testData5[3066];
@(posedge clk);
#1;data_in = testData5[3067];
@(posedge clk);
#1;data_in = testData5[3068];
@(posedge clk);
#1;data_in = testData5[3069];
@(posedge clk);
#1;data_in = testData5[3070];
@(posedge clk);
#1;data_in = testData5[3071];
@(posedge clk);
#1;data_in = testData5[3072];
@(posedge clk);
#1;data_in = testData5[3073];
@(posedge clk);
#1;data_in = testData5[3074];
@(posedge clk);
#1;data_in = testData5[3075];
@(posedge clk);
#1;data_in = testData5[3076];
@(posedge clk);
#1;data_in = testData5[3077];
@(posedge clk);
#1;data_in = testData5[3078];
@(posedge clk);
#1;data_in = testData5[3079];
@(posedge clk);
#1;data_in = testData5[3080];
@(posedge clk);
#1;data_in = testData5[3081];
@(posedge clk);
#1;data_in = testData5[3082];
@(posedge clk);
#1;data_in = testData5[3083];
@(posedge clk);
#1;data_in = testData5[3084];
@(posedge clk);
#1;data_in = testData5[3085];
@(posedge clk);
#1;data_in = testData5[3086];
@(posedge clk);
#1;data_in = testData5[3087];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3088]; 
@(posedge clk);
#1;data_in = testData5[3089];
@(posedge clk);
#1;data_in = testData5[3090];
@(posedge clk);
#1;data_in = testData5[3091];
@(posedge clk);
#1;data_in = testData5[3092];
@(posedge clk);
#1;data_in = testData5[3093];
@(posedge clk);
#1;data_in = testData5[3094];
@(posedge clk);
#1;data_in = testData5[3095];
@(posedge clk);
#1;data_in = testData5[3096];
@(posedge clk);
#1;data_in = testData5[3097];
@(posedge clk);
#1;data_in = testData5[3098];
@(posedge clk);
#1;data_in = testData5[3099];
@(posedge clk);
#1;data_in = testData5[3100];
@(posedge clk);
#1;data_in = testData5[3101];
@(posedge clk);
#1;data_in = testData5[3102];
@(posedge clk);
#1;data_in = testData5[3103];
@(posedge clk);
#1;data_in = testData5[3104];
@(posedge clk);
#1;data_in = testData5[3105];
@(posedge clk);
#1;data_in = testData5[3106];
@(posedge clk);
#1;data_in = testData5[3107];
@(posedge clk);
#1;data_in = testData5[3108];
@(posedge clk);
#1;data_in = testData5[3109];
@(posedge clk);
#1;data_in = testData5[3110];
@(posedge clk);
#1;data_in = testData5[3111];
@(posedge clk);
#1;data_in = testData5[3112];
@(posedge clk);
#1;data_in = testData5[3113];
@(posedge clk);
#1;data_in = testData5[3114];
@(posedge clk);
#1;data_in = testData5[3115];
@(posedge clk);
#1;data_in = testData5[3116];
@(posedge clk);
#1;data_in = testData5[3117];
@(posedge clk);
#1;data_in = testData5[3118];
@(posedge clk);
#1;data_in = testData5[3119];
@(posedge clk);
#1;data_in = testData5[3120];
@(posedge clk);
#1;data_in = testData5[3121];
@(posedge clk);
#1;data_in = testData5[3122];
@(posedge clk);
#1;data_in = testData5[3123];
@(posedge clk);
#1;data_in = testData5[3124];
@(posedge clk);
#1;data_in = testData5[3125];
@(posedge clk);
#1;data_in = testData5[3126];
@(posedge clk);
#1;data_in = testData5[3127];
@(posedge clk);
#1;data_in = testData5[3128];
@(posedge clk);
#1;data_in = testData5[3129];
@(posedge clk);
#1;data_in = testData5[3130];
@(posedge clk);
#1;data_in = testData5[3131];
@(posedge clk);
#1;data_in = testData5[3132];
@(posedge clk);
#1;data_in = testData5[3133];
@(posedge clk);
#1;data_in = testData5[3134];
@(posedge clk);
#1;data_in = testData5[3135];
@(posedge clk);
#1;data_in = testData5[3136];
@(posedge clk);
#1;data_in = testData5[3137];
@(posedge clk);
#1;data_in = testData5[3138];
@(posedge clk);
#1;data_in = testData5[3139];
@(posedge clk);
#1;data_in = testData5[3140];
@(posedge clk);
#1;data_in = testData5[3141];
@(posedge clk);
#1;data_in = testData5[3142];
@(posedge clk);
#1;data_in = testData5[3143];
@(posedge clk);
#1;data_in = testData5[3144];
@(posedge clk);
#1;data_in = testData5[3145];
@(posedge clk);
#1;data_in = testData5[3146];
@(posedge clk);
#1;data_in = testData5[3147];
@(posedge clk);
#1;data_in = testData5[3148];
@(posedge clk);
#1;data_in = testData5[3149];
@(posedge clk);
#1;data_in = testData5[3150];
@(posedge clk);
#1;data_in = testData5[3151];
@(posedge clk);
#1;data_in = testData5[3152];
@(posedge clk);
#1;data_in = testData5[3153];
@(posedge clk);
#1;data_in = testData5[3154];
@(posedge clk);
#1;data_in = testData5[3155];
@(posedge clk);
#1;data_in = testData5[3156];
@(posedge clk);
#1;data_in = testData5[3157];
@(posedge clk);
#1;data_in = testData5[3158];
@(posedge clk);
#1;data_in = testData5[3159];
@(posedge clk);
#1;data_in = testData5[3160];
@(posedge clk);
#1;data_in = testData5[3161];
@(posedge clk);
#1;data_in = testData5[3162];
@(posedge clk);
#1;data_in = testData5[3163];
@(posedge clk);
#1;data_in = testData5[3164];
@(posedge clk);
#1;data_in = testData5[3165];
@(posedge clk);
#1;data_in = testData5[3166];
@(posedge clk);
#1;data_in = testData5[3167];
@(posedge clk);
#1;data_in = testData5[3168];
@(posedge clk);
#1;data_in = testData5[3169];
@(posedge clk);
#1;data_in = testData5[3170];
@(posedge clk);
#1;data_in = testData5[3171];
@(posedge clk);
#1;data_in = testData5[3172];
@(posedge clk);
#1;data_in = testData5[3173];
@(posedge clk);
#1;data_in = testData5[3174];
@(posedge clk);
#1;data_in = testData5[3175];
@(posedge clk);
#1;data_in = testData5[3176];
@(posedge clk);
#1;data_in = testData5[3177];
@(posedge clk);
#1;data_in = testData5[3178];
@(posedge clk);
#1;data_in = testData5[3179];
@(posedge clk);
#1;data_in = testData5[3180];
@(posedge clk);
#1;data_in = testData5[3181];
@(posedge clk);
#1;data_in = testData5[3182];
@(posedge clk);
#1;data_in = testData5[3183];
@(posedge clk);
#1;data_in = testData5[3184];
@(posedge clk);
#1;data_in = testData5[3185];
@(posedge clk);
#1;data_in = testData5[3186];
@(posedge clk);
#1;data_in = testData5[3187];
@(posedge clk);
#1;data_in = testData5[3188];
@(posedge clk);
#1;data_in = testData5[3189];
@(posedge clk);
#1;data_in = testData5[3190];
@(posedge clk);
#1;data_in = testData5[3191];
@(posedge clk);
#1;data_in = testData5[3192];
@(posedge clk);
#1;data_in = testData5[3193];
@(posedge clk);
#1;data_in = testData5[3194];
@(posedge clk);
#1;data_in = testData5[3195];
@(posedge clk);
#1;data_in = testData5[3196];
@(posedge clk);
#1;data_in = testData5[3197];
@(posedge clk);
#1;data_in = testData5[3198];
@(posedge clk);
#1;data_in = testData5[3199];
@(posedge clk);
#1;data_in = testData5[3200];
@(posedge clk);
#1;data_in = testData5[3201];
@(posedge clk);
#1;data_in = testData5[3202];
@(posedge clk);
#1;data_in = testData5[3203];
@(posedge clk);
#1;data_in = testData5[3204];
@(posedge clk);
#1;data_in = testData5[3205];
@(posedge clk);
#1;data_in = testData5[3206];
@(posedge clk);
#1;data_in = testData5[3207];
@(posedge clk);
#1;data_in = testData5[3208];
@(posedge clk);
#1;data_in = testData5[3209];
@(posedge clk);
#1;data_in = testData5[3210];
@(posedge clk);
#1;data_in = testData5[3211];
@(posedge clk);
#1;data_in = testData5[3212];
@(posedge clk);
#1;data_in = testData5[3213];
@(posedge clk);
#1;data_in = testData5[3214];
@(posedge clk);
#1;data_in = testData5[3215];
@(posedge clk);
#1;data_in = testData5[3216];
@(posedge clk);
#1;data_in = testData5[3217];
@(posedge clk);
#1;data_in = testData5[3218];
@(posedge clk);
#1;data_in = testData5[3219];
@(posedge clk);
#1;data_in = testData5[3220];
@(posedge clk);
#1;data_in = testData5[3221];
@(posedge clk);
#1;data_in = testData5[3222];
@(posedge clk);
#1;data_in = testData5[3223];
@(posedge clk);
#1;data_in = testData5[3224];
@(posedge clk);
#1;data_in = testData5[3225];
@(posedge clk);
#1;data_in = testData5[3226];
@(posedge clk);
#1;data_in = testData5[3227];
@(posedge clk);
#1;data_in = testData5[3228];
@(posedge clk);
#1;data_in = testData5[3229];
@(posedge clk);
#1;data_in = testData5[3230];
@(posedge clk);
#1;data_in = testData5[3231];
@(posedge clk);
#1;data_in = testData5[3232];
@(posedge clk);
#1;data_in = testData5[3233];
@(posedge clk);
#1;data_in = testData5[3234];
@(posedge clk);
#1;data_in = testData5[3235];
@(posedge clk);
#1;data_in = testData5[3236];
@(posedge clk);
#1;data_in = testData5[3237];
@(posedge clk);
#1;data_in = testData5[3238];
@(posedge clk);
#1;data_in = testData5[3239];
@(posedge clk);
#1;data_in = testData5[3240];
@(posedge clk);
#1;data_in = testData5[3241];
@(posedge clk);
#1;data_in = testData5[3242];
@(posedge clk);
#1;data_in = testData5[3243];
@(posedge clk);
#1;data_in = testData5[3244];
@(posedge clk);
#1;data_in = testData5[3245];
@(posedge clk);
#1;data_in = testData5[3246];
@(posedge clk);
#1;data_in = testData5[3247];
@(posedge clk);
#1;data_in = testData5[3248];
@(posedge clk);
#1;data_in = testData5[3249];
@(posedge clk);
#1;data_in = testData5[3250];
@(posedge clk);
#1;data_in = testData5[3251];
@(posedge clk);
#1;data_in = testData5[3252];
@(posedge clk);
#1;data_in = testData5[3253];
@(posedge clk);
#1;data_in = testData5[3254];
@(posedge clk);
#1;data_in = testData5[3255];
@(posedge clk);
#1;data_in = testData5[3256];
@(posedge clk);
#1;data_in = testData5[3257];
@(posedge clk);
#1;data_in = testData5[3258];
@(posedge clk);
#1;data_in = testData5[3259];
@(posedge clk);
#1;data_in = testData5[3260];
@(posedge clk);
#1;data_in = testData5[3261];
@(posedge clk);
#1;data_in = testData5[3262];
@(posedge clk);
#1;data_in = testData5[3263];
@(posedge clk);
#1;data_in = testData5[3264];
@(posedge clk);
#1;data_in = testData5[3265];
@(posedge clk);
#1;data_in = testData5[3266];
@(posedge clk);
#1;data_in = testData5[3267];
@(posedge clk);
#1;data_in = testData5[3268];
@(posedge clk);
#1;data_in = testData5[3269];
@(posedge clk);
#1;data_in = testData5[3270];
@(posedge clk);
#1;data_in = testData5[3271];
@(posedge clk);
#1;data_in = testData5[3272];
@(posedge clk);
#1;data_in = testData5[3273];
@(posedge clk);
#1;data_in = testData5[3274];
@(posedge clk);
#1;data_in = testData5[3275];
@(posedge clk);
#1;data_in = testData5[3276];
@(posedge clk);
#1;data_in = testData5[3277];
@(posedge clk);
#1;data_in = testData5[3278];
@(posedge clk);
#1;data_in = testData5[3279];
@(posedge clk);
#1;data_in = testData5[3280];
@(posedge clk);
#1;data_in = testData5[3281];
@(posedge clk);
#1;data_in = testData5[3282];
@(posedge clk);
#1;data_in = testData5[3283];
@(posedge clk);
#1;data_in = testData5[3284];
@(posedge clk);
#1;data_in = testData5[3285];
@(posedge clk);
#1;data_in = testData5[3286];
@(posedge clk);
#1;data_in = testData5[3287];
@(posedge clk);
#1;data_in = testData5[3288];
@(posedge clk);
#1;data_in = testData5[3289];
@(posedge clk);
#1;data_in = testData5[3290];
@(posedge clk);
#1;data_in = testData5[3291];
@(posedge clk);
#1;data_in = testData5[3292];
@(posedge clk);
#1;data_in = testData5[3293];
@(posedge clk);
#1;data_in = testData5[3294];
@(posedge clk);
#1;data_in = testData5[3295];
@(posedge clk);
#1;data_in = testData5[3296];
@(posedge clk);
#1;data_in = testData5[3297];
@(posedge clk);
#1;data_in = testData5[3298];
@(posedge clk);
#1;data_in = testData5[3299];
@(posedge clk);
#1;data_in = testData5[3300];
@(posedge clk);
#1;data_in = testData5[3301];
@(posedge clk);
#1;data_in = testData5[3302];
@(posedge clk);
#1;data_in = testData5[3303];
@(posedge clk);
#1;data_in = testData5[3304];
@(posedge clk);
#1;data_in = testData5[3305];
@(posedge clk);
#1;data_in = testData5[3306];
@(posedge clk);
#1;data_in = testData5[3307];
@(posedge clk);
#1;data_in = testData5[3308];
@(posedge clk);
#1;data_in = testData5[3309];
@(posedge clk);
#1;data_in = testData5[3310];
@(posedge clk);
#1;data_in = testData5[3311];
@(posedge clk);
#1;data_in = testData5[3312];
@(posedge clk);
#1;data_in = testData5[3313];
@(posedge clk);
#1;data_in = testData5[3314];
@(posedge clk);
#1;data_in = testData5[3315];
@(posedge clk);
#1;data_in = testData5[3316];
@(posedge clk);
#1;data_in = testData5[3317];
@(posedge clk);
#1;data_in = testData5[3318];
@(posedge clk);
#1;data_in = testData5[3319];
@(posedge clk);
#1;data_in = testData5[3320];
@(posedge clk);
#1;data_in = testData5[3321];
@(posedge clk);
#1;data_in = testData5[3322];
@(posedge clk);
#1;data_in = testData5[3323];
@(posedge clk);
#1;data_in = testData5[3324];
@(posedge clk);
#1;data_in = testData5[3325];
@(posedge clk);
#1;data_in = testData5[3326];
@(posedge clk);
#1;data_in = testData5[3327];
@(posedge clk);
#1;data_in = testData5[3328];
@(posedge clk);
#1;data_in = testData5[3329];
@(posedge clk);
#1;data_in = testData5[3330];
@(posedge clk);
#1;data_in = testData5[3331];
@(posedge clk);
#1;data_in = testData5[3332];
@(posedge clk);
#1;data_in = testData5[3333];
@(posedge clk);
#1;data_in = testData5[3334];
@(posedge clk);
#1;data_in = testData5[3335];
@(posedge clk);
#1;data_in = testData5[3336];
@(posedge clk);
#1;data_in = testData5[3337];
@(posedge clk);
#1;data_in = testData5[3338];
@(posedge clk);
#1;data_in = testData5[3339];
@(posedge clk);
#1;data_in = testData5[3340];
@(posedge clk);
#1;data_in = testData5[3341];
@(posedge clk);
#1;data_in = testData5[3342];
@(posedge clk);
#1;data_in = testData5[3343];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3344]; 
@(posedge clk);
#1;data_in = testData5[3345];
@(posedge clk);
#1;data_in = testData5[3346];
@(posedge clk);
#1;data_in = testData5[3347];
@(posedge clk);
#1;data_in = testData5[3348];
@(posedge clk);
#1;data_in = testData5[3349];
@(posedge clk);
#1;data_in = testData5[3350];
@(posedge clk);
#1;data_in = testData5[3351];
@(posedge clk);
#1;data_in = testData5[3352];
@(posedge clk);
#1;data_in = testData5[3353];
@(posedge clk);
#1;data_in = testData5[3354];
@(posedge clk);
#1;data_in = testData5[3355];
@(posedge clk);
#1;data_in = testData5[3356];
@(posedge clk);
#1;data_in = testData5[3357];
@(posedge clk);
#1;data_in = testData5[3358];
@(posedge clk);
#1;data_in = testData5[3359];
@(posedge clk);
#1;data_in = testData5[3360];
@(posedge clk);
#1;data_in = testData5[3361];
@(posedge clk);
#1;data_in = testData5[3362];
@(posedge clk);
#1;data_in = testData5[3363];
@(posedge clk);
#1;data_in = testData5[3364];
@(posedge clk);
#1;data_in = testData5[3365];
@(posedge clk);
#1;data_in = testData5[3366];
@(posedge clk);
#1;data_in = testData5[3367];
@(posedge clk);
#1;data_in = testData5[3368];
@(posedge clk);
#1;data_in = testData5[3369];
@(posedge clk);
#1;data_in = testData5[3370];
@(posedge clk);
#1;data_in = testData5[3371];
@(posedge clk);
#1;data_in = testData5[3372];
@(posedge clk);
#1;data_in = testData5[3373];
@(posedge clk);
#1;data_in = testData5[3374];
@(posedge clk);
#1;data_in = testData5[3375];
@(posedge clk);
#1;data_in = testData5[3376];
@(posedge clk);
#1;data_in = testData5[3377];
@(posedge clk);
#1;data_in = testData5[3378];
@(posedge clk);
#1;data_in = testData5[3379];
@(posedge clk);
#1;data_in = testData5[3380];
@(posedge clk);
#1;data_in = testData5[3381];
@(posedge clk);
#1;data_in = testData5[3382];
@(posedge clk);
#1;data_in = testData5[3383];
@(posedge clk);
#1;data_in = testData5[3384];
@(posedge clk);
#1;data_in = testData5[3385];
@(posedge clk);
#1;data_in = testData5[3386];
@(posedge clk);
#1;data_in = testData5[3387];
@(posedge clk);
#1;data_in = testData5[3388];
@(posedge clk);
#1;data_in = testData5[3389];
@(posedge clk);
#1;data_in = testData5[3390];
@(posedge clk);
#1;data_in = testData5[3391];
@(posedge clk);
#1;data_in = testData5[3392];
@(posedge clk);
#1;data_in = testData5[3393];
@(posedge clk);
#1;data_in = testData5[3394];
@(posedge clk);
#1;data_in = testData5[3395];
@(posedge clk);
#1;data_in = testData5[3396];
@(posedge clk);
#1;data_in = testData5[3397];
@(posedge clk);
#1;data_in = testData5[3398];
@(posedge clk);
#1;data_in = testData5[3399];
@(posedge clk);
#1;data_in = testData5[3400];
@(posedge clk);
#1;data_in = testData5[3401];
@(posedge clk);
#1;data_in = testData5[3402];
@(posedge clk);
#1;data_in = testData5[3403];
@(posedge clk);
#1;data_in = testData5[3404];
@(posedge clk);
#1;data_in = testData5[3405];
@(posedge clk);
#1;data_in = testData5[3406];
@(posedge clk);
#1;data_in = testData5[3407];
@(posedge clk);
#1;data_in = testData5[3408];
@(posedge clk);
#1;data_in = testData5[3409];
@(posedge clk);
#1;data_in = testData5[3410];
@(posedge clk);
#1;data_in = testData5[3411];
@(posedge clk);
#1;data_in = testData5[3412];
@(posedge clk);
#1;data_in = testData5[3413];
@(posedge clk);
#1;data_in = testData5[3414];
@(posedge clk);
#1;data_in = testData5[3415];
@(posedge clk);
#1;data_in = testData5[3416];
@(posedge clk);
#1;data_in = testData5[3417];
@(posedge clk);
#1;data_in = testData5[3418];
@(posedge clk);
#1;data_in = testData5[3419];
@(posedge clk);
#1;data_in = testData5[3420];
@(posedge clk);
#1;data_in = testData5[3421];
@(posedge clk);
#1;data_in = testData5[3422];
@(posedge clk);
#1;data_in = testData5[3423];
@(posedge clk);
#1;data_in = testData5[3424];
@(posedge clk);
#1;data_in = testData5[3425];
@(posedge clk);
#1;data_in = testData5[3426];
@(posedge clk);
#1;data_in = testData5[3427];
@(posedge clk);
#1;data_in = testData5[3428];
@(posedge clk);
#1;data_in = testData5[3429];
@(posedge clk);
#1;data_in = testData5[3430];
@(posedge clk);
#1;data_in = testData5[3431];
@(posedge clk);
#1;data_in = testData5[3432];
@(posedge clk);
#1;data_in = testData5[3433];
@(posedge clk);
#1;data_in = testData5[3434];
@(posedge clk);
#1;data_in = testData5[3435];
@(posedge clk);
#1;data_in = testData5[3436];
@(posedge clk);
#1;data_in = testData5[3437];
@(posedge clk);
#1;data_in = testData5[3438];
@(posedge clk);
#1;data_in = testData5[3439];
@(posedge clk);
#1;data_in = testData5[3440];
@(posedge clk);
#1;data_in = testData5[3441];
@(posedge clk);
#1;data_in = testData5[3442];
@(posedge clk);
#1;data_in = testData5[3443];
@(posedge clk);
#1;data_in = testData5[3444];
@(posedge clk);
#1;data_in = testData5[3445];
@(posedge clk);
#1;data_in = testData5[3446];
@(posedge clk);
#1;data_in = testData5[3447];
@(posedge clk);
#1;data_in = testData5[3448];
@(posedge clk);
#1;data_in = testData5[3449];
@(posedge clk);
#1;data_in = testData5[3450];
@(posedge clk);
#1;data_in = testData5[3451];
@(posedge clk);
#1;data_in = testData5[3452];
@(posedge clk);
#1;data_in = testData5[3453];
@(posedge clk);
#1;data_in = testData5[3454];
@(posedge clk);
#1;data_in = testData5[3455];
@(posedge clk);
#1;data_in = testData5[3456];
@(posedge clk);
#1;data_in = testData5[3457];
@(posedge clk);
#1;data_in = testData5[3458];
@(posedge clk);
#1;data_in = testData5[3459];
@(posedge clk);
#1;data_in = testData5[3460];
@(posedge clk);
#1;data_in = testData5[3461];
@(posedge clk);
#1;data_in = testData5[3462];
@(posedge clk);
#1;data_in = testData5[3463];
@(posedge clk);
#1;data_in = testData5[3464];
@(posedge clk);
#1;data_in = testData5[3465];
@(posedge clk);
#1;data_in = testData5[3466];
@(posedge clk);
#1;data_in = testData5[3467];
@(posedge clk);
#1;data_in = testData5[3468];
@(posedge clk);
#1;data_in = testData5[3469];
@(posedge clk);
#1;data_in = testData5[3470];
@(posedge clk);
#1;data_in = testData5[3471];
@(posedge clk);
#1;data_in = testData5[3472];
@(posedge clk);
#1;data_in = testData5[3473];
@(posedge clk);
#1;data_in = testData5[3474];
@(posedge clk);
#1;data_in = testData5[3475];
@(posedge clk);
#1;data_in = testData5[3476];
@(posedge clk);
#1;data_in = testData5[3477];
@(posedge clk);
#1;data_in = testData5[3478];
@(posedge clk);
#1;data_in = testData5[3479];
@(posedge clk);
#1;data_in = testData5[3480];
@(posedge clk);
#1;data_in = testData5[3481];
@(posedge clk);
#1;data_in = testData5[3482];
@(posedge clk);
#1;data_in = testData5[3483];
@(posedge clk);
#1;data_in = testData5[3484];
@(posedge clk);
#1;data_in = testData5[3485];
@(posedge clk);
#1;data_in = testData5[3486];
@(posedge clk);
#1;data_in = testData5[3487];
@(posedge clk);
#1;data_in = testData5[3488];
@(posedge clk);
#1;data_in = testData5[3489];
@(posedge clk);
#1;data_in = testData5[3490];
@(posedge clk);
#1;data_in = testData5[3491];
@(posedge clk);
#1;data_in = testData5[3492];
@(posedge clk);
#1;data_in = testData5[3493];
@(posedge clk);
#1;data_in = testData5[3494];
@(posedge clk);
#1;data_in = testData5[3495];
@(posedge clk);
#1;data_in = testData5[3496];
@(posedge clk);
#1;data_in = testData5[3497];
@(posedge clk);
#1;data_in = testData5[3498];
@(posedge clk);
#1;data_in = testData5[3499];
@(posedge clk);
#1;data_in = testData5[3500];
@(posedge clk);
#1;data_in = testData5[3501];
@(posedge clk);
#1;data_in = testData5[3502];
@(posedge clk);
#1;data_in = testData5[3503];
@(posedge clk);
#1;data_in = testData5[3504];
@(posedge clk);
#1;data_in = testData5[3505];
@(posedge clk);
#1;data_in = testData5[3506];
@(posedge clk);
#1;data_in = testData5[3507];
@(posedge clk);
#1;data_in = testData5[3508];
@(posedge clk);
#1;data_in = testData5[3509];
@(posedge clk);
#1;data_in = testData5[3510];
@(posedge clk);
#1;data_in = testData5[3511];
@(posedge clk);
#1;data_in = testData5[3512];
@(posedge clk);
#1;data_in = testData5[3513];
@(posedge clk);
#1;data_in = testData5[3514];
@(posedge clk);
#1;data_in = testData5[3515];
@(posedge clk);
#1;data_in = testData5[3516];
@(posedge clk);
#1;data_in = testData5[3517];
@(posedge clk);
#1;data_in = testData5[3518];
@(posedge clk);
#1;data_in = testData5[3519];
@(posedge clk);
#1;data_in = testData5[3520];
@(posedge clk);
#1;data_in = testData5[3521];
@(posedge clk);
#1;data_in = testData5[3522];
@(posedge clk);
#1;data_in = testData5[3523];
@(posedge clk);
#1;data_in = testData5[3524];
@(posedge clk);
#1;data_in = testData5[3525];
@(posedge clk);
#1;data_in = testData5[3526];
@(posedge clk);
#1;data_in = testData5[3527];
@(posedge clk);
#1;data_in = testData5[3528];
@(posedge clk);
#1;data_in = testData5[3529];
@(posedge clk);
#1;data_in = testData5[3530];
@(posedge clk);
#1;data_in = testData5[3531];
@(posedge clk);
#1;data_in = testData5[3532];
@(posedge clk);
#1;data_in = testData5[3533];
@(posedge clk);
#1;data_in = testData5[3534];
@(posedge clk);
#1;data_in = testData5[3535];
@(posedge clk);
#1;data_in = testData5[3536];
@(posedge clk);
#1;data_in = testData5[3537];
@(posedge clk);
#1;data_in = testData5[3538];
@(posedge clk);
#1;data_in = testData5[3539];
@(posedge clk);
#1;data_in = testData5[3540];
@(posedge clk);
#1;data_in = testData5[3541];
@(posedge clk);
#1;data_in = testData5[3542];
@(posedge clk);
#1;data_in = testData5[3543];
@(posedge clk);
#1;data_in = testData5[3544];
@(posedge clk);
#1;data_in = testData5[3545];
@(posedge clk);
#1;data_in = testData5[3546];
@(posedge clk);
#1;data_in = testData5[3547];
@(posedge clk);
#1;data_in = testData5[3548];
@(posedge clk);
#1;data_in = testData5[3549];
@(posedge clk);
#1;data_in = testData5[3550];
@(posedge clk);
#1;data_in = testData5[3551];
@(posedge clk);
#1;data_in = testData5[3552];
@(posedge clk);
#1;data_in = testData5[3553];
@(posedge clk);
#1;data_in = testData5[3554];
@(posedge clk);
#1;data_in = testData5[3555];
@(posedge clk);
#1;data_in = testData5[3556];
@(posedge clk);
#1;data_in = testData5[3557];
@(posedge clk);
#1;data_in = testData5[3558];
@(posedge clk);
#1;data_in = testData5[3559];
@(posedge clk);
#1;data_in = testData5[3560];
@(posedge clk);
#1;data_in = testData5[3561];
@(posedge clk);
#1;data_in = testData5[3562];
@(posedge clk);
#1;data_in = testData5[3563];
@(posedge clk);
#1;data_in = testData5[3564];
@(posedge clk);
#1;data_in = testData5[3565];
@(posedge clk);
#1;data_in = testData5[3566];
@(posedge clk);
#1;data_in = testData5[3567];
@(posedge clk);
#1;data_in = testData5[3568];
@(posedge clk);
#1;data_in = testData5[3569];
@(posedge clk);
#1;data_in = testData5[3570];
@(posedge clk);
#1;data_in = testData5[3571];
@(posedge clk);
#1;data_in = testData5[3572];
@(posedge clk);
#1;data_in = testData5[3573];
@(posedge clk);
#1;data_in = testData5[3574];
@(posedge clk);
#1;data_in = testData5[3575];
@(posedge clk);
#1;data_in = testData5[3576];
@(posedge clk);
#1;data_in = testData5[3577];
@(posedge clk);
#1;data_in = testData5[3578];
@(posedge clk);
#1;data_in = testData5[3579];
@(posedge clk);
#1;data_in = testData5[3580];
@(posedge clk);
#1;data_in = testData5[3581];
@(posedge clk);
#1;data_in = testData5[3582];
@(posedge clk);
#1;data_in = testData5[3583];
@(posedge clk);
#1;data_in = testData5[3584];
@(posedge clk);
#1;data_in = testData5[3585];
@(posedge clk);
#1;data_in = testData5[3586];
@(posedge clk);
#1;data_in = testData5[3587];
@(posedge clk);
#1;data_in = testData5[3588];
@(posedge clk);
#1;data_in = testData5[3589];
@(posedge clk);
#1;data_in = testData5[3590];
@(posedge clk);
#1;data_in = testData5[3591];
@(posedge clk);
#1;data_in = testData5[3592];
@(posedge clk);
#1;data_in = testData5[3593];
@(posedge clk);
#1;data_in = testData5[3594];
@(posedge clk);
#1;data_in = testData5[3595];
@(posedge clk);
#1;data_in = testData5[3596];
@(posedge clk);
#1;data_in = testData5[3597];
@(posedge clk);
#1;data_in = testData5[3598];
@(posedge clk);
#1;data_in = testData5[3599];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3600]; 
@(posedge clk);
#1;data_in = testData5[3601];
@(posedge clk);
#1;data_in = testData5[3602];
@(posedge clk);
#1;data_in = testData5[3603];
@(posedge clk);
#1;data_in = testData5[3604];
@(posedge clk);
#1;data_in = testData5[3605];
@(posedge clk);
#1;data_in = testData5[3606];
@(posedge clk);
#1;data_in = testData5[3607];
@(posedge clk);
#1;data_in = testData5[3608];
@(posedge clk);
#1;data_in = testData5[3609];
@(posedge clk);
#1;data_in = testData5[3610];
@(posedge clk);
#1;data_in = testData5[3611];
@(posedge clk);
#1;data_in = testData5[3612];
@(posedge clk);
#1;data_in = testData5[3613];
@(posedge clk);
#1;data_in = testData5[3614];
@(posedge clk);
#1;data_in = testData5[3615];
@(posedge clk);
#1;data_in = testData5[3616];
@(posedge clk);
#1;data_in = testData5[3617];
@(posedge clk);
#1;data_in = testData5[3618];
@(posedge clk);
#1;data_in = testData5[3619];
@(posedge clk);
#1;data_in = testData5[3620];
@(posedge clk);
#1;data_in = testData5[3621];
@(posedge clk);
#1;data_in = testData5[3622];
@(posedge clk);
#1;data_in = testData5[3623];
@(posedge clk);
#1;data_in = testData5[3624];
@(posedge clk);
#1;data_in = testData5[3625];
@(posedge clk);
#1;data_in = testData5[3626];
@(posedge clk);
#1;data_in = testData5[3627];
@(posedge clk);
#1;data_in = testData5[3628];
@(posedge clk);
#1;data_in = testData5[3629];
@(posedge clk);
#1;data_in = testData5[3630];
@(posedge clk);
#1;data_in = testData5[3631];
@(posedge clk);
#1;data_in = testData5[3632];
@(posedge clk);
#1;data_in = testData5[3633];
@(posedge clk);
#1;data_in = testData5[3634];
@(posedge clk);
#1;data_in = testData5[3635];
@(posedge clk);
#1;data_in = testData5[3636];
@(posedge clk);
#1;data_in = testData5[3637];
@(posedge clk);
#1;data_in = testData5[3638];
@(posedge clk);
#1;data_in = testData5[3639];
@(posedge clk);
#1;data_in = testData5[3640];
@(posedge clk);
#1;data_in = testData5[3641];
@(posedge clk);
#1;data_in = testData5[3642];
@(posedge clk);
#1;data_in = testData5[3643];
@(posedge clk);
#1;data_in = testData5[3644];
@(posedge clk);
#1;data_in = testData5[3645];
@(posedge clk);
#1;data_in = testData5[3646];
@(posedge clk);
#1;data_in = testData5[3647];
@(posedge clk);
#1;data_in = testData5[3648];
@(posedge clk);
#1;data_in = testData5[3649];
@(posedge clk);
#1;data_in = testData5[3650];
@(posedge clk);
#1;data_in = testData5[3651];
@(posedge clk);
#1;data_in = testData5[3652];
@(posedge clk);
#1;data_in = testData5[3653];
@(posedge clk);
#1;data_in = testData5[3654];
@(posedge clk);
#1;data_in = testData5[3655];
@(posedge clk);
#1;data_in = testData5[3656];
@(posedge clk);
#1;data_in = testData5[3657];
@(posedge clk);
#1;data_in = testData5[3658];
@(posedge clk);
#1;data_in = testData5[3659];
@(posedge clk);
#1;data_in = testData5[3660];
@(posedge clk);
#1;data_in = testData5[3661];
@(posedge clk);
#1;data_in = testData5[3662];
@(posedge clk);
#1;data_in = testData5[3663];
@(posedge clk);
#1;data_in = testData5[3664];
@(posedge clk);
#1;data_in = testData5[3665];
@(posedge clk);
#1;data_in = testData5[3666];
@(posedge clk);
#1;data_in = testData5[3667];
@(posedge clk);
#1;data_in = testData5[3668];
@(posedge clk);
#1;data_in = testData5[3669];
@(posedge clk);
#1;data_in = testData5[3670];
@(posedge clk);
#1;data_in = testData5[3671];
@(posedge clk);
#1;data_in = testData5[3672];
@(posedge clk);
#1;data_in = testData5[3673];
@(posedge clk);
#1;data_in = testData5[3674];
@(posedge clk);
#1;data_in = testData5[3675];
@(posedge clk);
#1;data_in = testData5[3676];
@(posedge clk);
#1;data_in = testData5[3677];
@(posedge clk);
#1;data_in = testData5[3678];
@(posedge clk);
#1;data_in = testData5[3679];
@(posedge clk);
#1;data_in = testData5[3680];
@(posedge clk);
#1;data_in = testData5[3681];
@(posedge clk);
#1;data_in = testData5[3682];
@(posedge clk);
#1;data_in = testData5[3683];
@(posedge clk);
#1;data_in = testData5[3684];
@(posedge clk);
#1;data_in = testData5[3685];
@(posedge clk);
#1;data_in = testData5[3686];
@(posedge clk);
#1;data_in = testData5[3687];
@(posedge clk);
#1;data_in = testData5[3688];
@(posedge clk);
#1;data_in = testData5[3689];
@(posedge clk);
#1;data_in = testData5[3690];
@(posedge clk);
#1;data_in = testData5[3691];
@(posedge clk);
#1;data_in = testData5[3692];
@(posedge clk);
#1;data_in = testData5[3693];
@(posedge clk);
#1;data_in = testData5[3694];
@(posedge clk);
#1;data_in = testData5[3695];
@(posedge clk);
#1;data_in = testData5[3696];
@(posedge clk);
#1;data_in = testData5[3697];
@(posedge clk);
#1;data_in = testData5[3698];
@(posedge clk);
#1;data_in = testData5[3699];
@(posedge clk);
#1;data_in = testData5[3700];
@(posedge clk);
#1;data_in = testData5[3701];
@(posedge clk);
#1;data_in = testData5[3702];
@(posedge clk);
#1;data_in = testData5[3703];
@(posedge clk);
#1;data_in = testData5[3704];
@(posedge clk);
#1;data_in = testData5[3705];
@(posedge clk);
#1;data_in = testData5[3706];
@(posedge clk);
#1;data_in = testData5[3707];
@(posedge clk);
#1;data_in = testData5[3708];
@(posedge clk);
#1;data_in = testData5[3709];
@(posedge clk);
#1;data_in = testData5[3710];
@(posedge clk);
#1;data_in = testData5[3711];
@(posedge clk);
#1;data_in = testData5[3712];
@(posedge clk);
#1;data_in = testData5[3713];
@(posedge clk);
#1;data_in = testData5[3714];
@(posedge clk);
#1;data_in = testData5[3715];
@(posedge clk);
#1;data_in = testData5[3716];
@(posedge clk);
#1;data_in = testData5[3717];
@(posedge clk);
#1;data_in = testData5[3718];
@(posedge clk);
#1;data_in = testData5[3719];
@(posedge clk);
#1;data_in = testData5[3720];
@(posedge clk);
#1;data_in = testData5[3721];
@(posedge clk);
#1;data_in = testData5[3722];
@(posedge clk);
#1;data_in = testData5[3723];
@(posedge clk);
#1;data_in = testData5[3724];
@(posedge clk);
#1;data_in = testData5[3725];
@(posedge clk);
#1;data_in = testData5[3726];
@(posedge clk);
#1;data_in = testData5[3727];
@(posedge clk);
#1;data_in = testData5[3728];
@(posedge clk);
#1;data_in = testData5[3729];
@(posedge clk);
#1;data_in = testData5[3730];
@(posedge clk);
#1;data_in = testData5[3731];
@(posedge clk);
#1;data_in = testData5[3732];
@(posedge clk);
#1;data_in = testData5[3733];
@(posedge clk);
#1;data_in = testData5[3734];
@(posedge clk);
#1;data_in = testData5[3735];
@(posedge clk);
#1;data_in = testData5[3736];
@(posedge clk);
#1;data_in = testData5[3737];
@(posedge clk);
#1;data_in = testData5[3738];
@(posedge clk);
#1;data_in = testData5[3739];
@(posedge clk);
#1;data_in = testData5[3740];
@(posedge clk);
#1;data_in = testData5[3741];
@(posedge clk);
#1;data_in = testData5[3742];
@(posedge clk);
#1;data_in = testData5[3743];
@(posedge clk);
#1;data_in = testData5[3744];
@(posedge clk);
#1;data_in = testData5[3745];
@(posedge clk);
#1;data_in = testData5[3746];
@(posedge clk);
#1;data_in = testData5[3747];
@(posedge clk);
#1;data_in = testData5[3748];
@(posedge clk);
#1;data_in = testData5[3749];
@(posedge clk);
#1;data_in = testData5[3750];
@(posedge clk);
#1;data_in = testData5[3751];
@(posedge clk);
#1;data_in = testData5[3752];
@(posedge clk);
#1;data_in = testData5[3753];
@(posedge clk);
#1;data_in = testData5[3754];
@(posedge clk);
#1;data_in = testData5[3755];
@(posedge clk);
#1;data_in = testData5[3756];
@(posedge clk);
#1;data_in = testData5[3757];
@(posedge clk);
#1;data_in = testData5[3758];
@(posedge clk);
#1;data_in = testData5[3759];
@(posedge clk);
#1;data_in = testData5[3760];
@(posedge clk);
#1;data_in = testData5[3761];
@(posedge clk);
#1;data_in = testData5[3762];
@(posedge clk);
#1;data_in = testData5[3763];
@(posedge clk);
#1;data_in = testData5[3764];
@(posedge clk);
#1;data_in = testData5[3765];
@(posedge clk);
#1;data_in = testData5[3766];
@(posedge clk);
#1;data_in = testData5[3767];
@(posedge clk);
#1;data_in = testData5[3768];
@(posedge clk);
#1;data_in = testData5[3769];
@(posedge clk);
#1;data_in = testData5[3770];
@(posedge clk);
#1;data_in = testData5[3771];
@(posedge clk);
#1;data_in = testData5[3772];
@(posedge clk);
#1;data_in = testData5[3773];
@(posedge clk);
#1;data_in = testData5[3774];
@(posedge clk);
#1;data_in = testData5[3775];
@(posedge clk);
#1;data_in = testData5[3776];
@(posedge clk);
#1;data_in = testData5[3777];
@(posedge clk);
#1;data_in = testData5[3778];
@(posedge clk);
#1;data_in = testData5[3779];
@(posedge clk);
#1;data_in = testData5[3780];
@(posedge clk);
#1;data_in = testData5[3781];
@(posedge clk);
#1;data_in = testData5[3782];
@(posedge clk);
#1;data_in = testData5[3783];
@(posedge clk);
#1;data_in = testData5[3784];
@(posedge clk);
#1;data_in = testData5[3785];
@(posedge clk);
#1;data_in = testData5[3786];
@(posedge clk);
#1;data_in = testData5[3787];
@(posedge clk);
#1;data_in = testData5[3788];
@(posedge clk);
#1;data_in = testData5[3789];
@(posedge clk);
#1;data_in = testData5[3790];
@(posedge clk);
#1;data_in = testData5[3791];
@(posedge clk);
#1;data_in = testData5[3792];
@(posedge clk);
#1;data_in = testData5[3793];
@(posedge clk);
#1;data_in = testData5[3794];
@(posedge clk);
#1;data_in = testData5[3795];
@(posedge clk);
#1;data_in = testData5[3796];
@(posedge clk);
#1;data_in = testData5[3797];
@(posedge clk);
#1;data_in = testData5[3798];
@(posedge clk);
#1;data_in = testData5[3799];
@(posedge clk);
#1;data_in = testData5[3800];
@(posedge clk);
#1;data_in = testData5[3801];
@(posedge clk);
#1;data_in = testData5[3802];
@(posedge clk);
#1;data_in = testData5[3803];
@(posedge clk);
#1;data_in = testData5[3804];
@(posedge clk);
#1;data_in = testData5[3805];
@(posedge clk);
#1;data_in = testData5[3806];
@(posedge clk);
#1;data_in = testData5[3807];
@(posedge clk);
#1;data_in = testData5[3808];
@(posedge clk);
#1;data_in = testData5[3809];
@(posedge clk);
#1;data_in = testData5[3810];
@(posedge clk);
#1;data_in = testData5[3811];
@(posedge clk);
#1;data_in = testData5[3812];
@(posedge clk);
#1;data_in = testData5[3813];
@(posedge clk);
#1;data_in = testData5[3814];
@(posedge clk);
#1;data_in = testData5[3815];
@(posedge clk);
#1;data_in = testData5[3816];
@(posedge clk);
#1;data_in = testData5[3817];
@(posedge clk);
#1;data_in = testData5[3818];
@(posedge clk);
#1;data_in = testData5[3819];
@(posedge clk);
#1;data_in = testData5[3820];
@(posedge clk);
#1;data_in = testData5[3821];
@(posedge clk);
#1;data_in = testData5[3822];
@(posedge clk);
#1;data_in = testData5[3823];
@(posedge clk);
#1;data_in = testData5[3824];
@(posedge clk);
#1;data_in = testData5[3825];
@(posedge clk);
#1;data_in = testData5[3826];
@(posedge clk);
#1;data_in = testData5[3827];
@(posedge clk);
#1;data_in = testData5[3828];
@(posedge clk);
#1;data_in = testData5[3829];
@(posedge clk);
#1;data_in = testData5[3830];
@(posedge clk);
#1;data_in = testData5[3831];
@(posedge clk);
#1;data_in = testData5[3832];
@(posedge clk);
#1;data_in = testData5[3833];
@(posedge clk);
#1;data_in = testData5[3834];
@(posedge clk);
#1;data_in = testData5[3835];
@(posedge clk);
#1;data_in = testData5[3836];
@(posedge clk);
#1;data_in = testData5[3837];
@(posedge clk);
#1;data_in = testData5[3838];
@(posedge clk);
#1;data_in = testData5[3839];
@(posedge clk);
#1;data_in = testData5[3840];
@(posedge clk);
#1;data_in = testData5[3841];
@(posedge clk);
#1;data_in = testData5[3842];
@(posedge clk);
#1;data_in = testData5[3843];
@(posedge clk);
#1;data_in = testData5[3844];
@(posedge clk);
#1;data_in = testData5[3845];
@(posedge clk);
#1;data_in = testData5[3846];
@(posedge clk);
#1;data_in = testData5[3847];
@(posedge clk);
#1;data_in = testData5[3848];
@(posedge clk);
#1;data_in = testData5[3849];
@(posedge clk);
#1;data_in = testData5[3850];
@(posedge clk);
#1;data_in = testData5[3851];
@(posedge clk);
#1;data_in = testData5[3852];
@(posedge clk);
#1;data_in = testData5[3853];
@(posedge clk);
#1;data_in = testData5[3854];
@(posedge clk);
#1;data_in = testData5[3855];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3856]; 
@(posedge clk);
#1;data_in = testData5[3857];
@(posedge clk);
#1;data_in = testData5[3858];
@(posedge clk);
#1;data_in = testData5[3859];
@(posedge clk);
#1;data_in = testData5[3860];
@(posedge clk);
#1;data_in = testData5[3861];
@(posedge clk);
#1;data_in = testData5[3862];
@(posedge clk);
#1;data_in = testData5[3863];
@(posedge clk);
#1;data_in = testData5[3864];
@(posedge clk);
#1;data_in = testData5[3865];
@(posedge clk);
#1;data_in = testData5[3866];
@(posedge clk);
#1;data_in = testData5[3867];
@(posedge clk);
#1;data_in = testData5[3868];
@(posedge clk);
#1;data_in = testData5[3869];
@(posedge clk);
#1;data_in = testData5[3870];
@(posedge clk);
#1;data_in = testData5[3871];
@(posedge clk);
#1;data_in = testData5[3872];
@(posedge clk);
#1;data_in = testData5[3873];
@(posedge clk);
#1;data_in = testData5[3874];
@(posedge clk);
#1;data_in = testData5[3875];
@(posedge clk);
#1;data_in = testData5[3876];
@(posedge clk);
#1;data_in = testData5[3877];
@(posedge clk);
#1;data_in = testData5[3878];
@(posedge clk);
#1;data_in = testData5[3879];
@(posedge clk);
#1;data_in = testData5[3880];
@(posedge clk);
#1;data_in = testData5[3881];
@(posedge clk);
#1;data_in = testData5[3882];
@(posedge clk);
#1;data_in = testData5[3883];
@(posedge clk);
#1;data_in = testData5[3884];
@(posedge clk);
#1;data_in = testData5[3885];
@(posedge clk);
#1;data_in = testData5[3886];
@(posedge clk);
#1;data_in = testData5[3887];
@(posedge clk);
#1;data_in = testData5[3888];
@(posedge clk);
#1;data_in = testData5[3889];
@(posedge clk);
#1;data_in = testData5[3890];
@(posedge clk);
#1;data_in = testData5[3891];
@(posedge clk);
#1;data_in = testData5[3892];
@(posedge clk);
#1;data_in = testData5[3893];
@(posedge clk);
#1;data_in = testData5[3894];
@(posedge clk);
#1;data_in = testData5[3895];
@(posedge clk);
#1;data_in = testData5[3896];
@(posedge clk);
#1;data_in = testData5[3897];
@(posedge clk);
#1;data_in = testData5[3898];
@(posedge clk);
#1;data_in = testData5[3899];
@(posedge clk);
#1;data_in = testData5[3900];
@(posedge clk);
#1;data_in = testData5[3901];
@(posedge clk);
#1;data_in = testData5[3902];
@(posedge clk);
#1;data_in = testData5[3903];
@(posedge clk);
#1;data_in = testData5[3904];
@(posedge clk);
#1;data_in = testData5[3905];
@(posedge clk);
#1;data_in = testData5[3906];
@(posedge clk);
#1;data_in = testData5[3907];
@(posedge clk);
#1;data_in = testData5[3908];
@(posedge clk);
#1;data_in = testData5[3909];
@(posedge clk);
#1;data_in = testData5[3910];
@(posedge clk);
#1;data_in = testData5[3911];
@(posedge clk);
#1;data_in = testData5[3912];
@(posedge clk);
#1;data_in = testData5[3913];
@(posedge clk);
#1;data_in = testData5[3914];
@(posedge clk);
#1;data_in = testData5[3915];
@(posedge clk);
#1;data_in = testData5[3916];
@(posedge clk);
#1;data_in = testData5[3917];
@(posedge clk);
#1;data_in = testData5[3918];
@(posedge clk);
#1;data_in = testData5[3919];
@(posedge clk);
#1;data_in = testData5[3920];
@(posedge clk);
#1;data_in = testData5[3921];
@(posedge clk);
#1;data_in = testData5[3922];
@(posedge clk);
#1;data_in = testData5[3923];
@(posedge clk);
#1;data_in = testData5[3924];
@(posedge clk);
#1;data_in = testData5[3925];
@(posedge clk);
#1;data_in = testData5[3926];
@(posedge clk);
#1;data_in = testData5[3927];
@(posedge clk);
#1;data_in = testData5[3928];
@(posedge clk);
#1;data_in = testData5[3929];
@(posedge clk);
#1;data_in = testData5[3930];
@(posedge clk);
#1;data_in = testData5[3931];
@(posedge clk);
#1;data_in = testData5[3932];
@(posedge clk);
#1;data_in = testData5[3933];
@(posedge clk);
#1;data_in = testData5[3934];
@(posedge clk);
#1;data_in = testData5[3935];
@(posedge clk);
#1;data_in = testData5[3936];
@(posedge clk);
#1;data_in = testData5[3937];
@(posedge clk);
#1;data_in = testData5[3938];
@(posedge clk);
#1;data_in = testData5[3939];
@(posedge clk);
#1;data_in = testData5[3940];
@(posedge clk);
#1;data_in = testData5[3941];
@(posedge clk);
#1;data_in = testData5[3942];
@(posedge clk);
#1;data_in = testData5[3943];
@(posedge clk);
#1;data_in = testData5[3944];
@(posedge clk);
#1;data_in = testData5[3945];
@(posedge clk);
#1;data_in = testData5[3946];
@(posedge clk);
#1;data_in = testData5[3947];
@(posedge clk);
#1;data_in = testData5[3948];
@(posedge clk);
#1;data_in = testData5[3949];
@(posedge clk);
#1;data_in = testData5[3950];
@(posedge clk);
#1;data_in = testData5[3951];
@(posedge clk);
#1;data_in = testData5[3952];
@(posedge clk);
#1;data_in = testData5[3953];
@(posedge clk);
#1;data_in = testData5[3954];
@(posedge clk);
#1;data_in = testData5[3955];
@(posedge clk);
#1;data_in = testData5[3956];
@(posedge clk);
#1;data_in = testData5[3957];
@(posedge clk);
#1;data_in = testData5[3958];
@(posedge clk);
#1;data_in = testData5[3959];
@(posedge clk);
#1;data_in = testData5[3960];
@(posedge clk);
#1;data_in = testData5[3961];
@(posedge clk);
#1;data_in = testData5[3962];
@(posedge clk);
#1;data_in = testData5[3963];
@(posedge clk);
#1;data_in = testData5[3964];
@(posedge clk);
#1;data_in = testData5[3965];
@(posedge clk);
#1;data_in = testData5[3966];
@(posedge clk);
#1;data_in = testData5[3967];
@(posedge clk);
#1;data_in = testData5[3968];
@(posedge clk);
#1;data_in = testData5[3969];
@(posedge clk);
#1;data_in = testData5[3970];
@(posedge clk);
#1;data_in = testData5[3971];
@(posedge clk);
#1;data_in = testData5[3972];
@(posedge clk);
#1;data_in = testData5[3973];
@(posedge clk);
#1;data_in = testData5[3974];
@(posedge clk);
#1;data_in = testData5[3975];
@(posedge clk);
#1;data_in = testData5[3976];
@(posedge clk);
#1;data_in = testData5[3977];
@(posedge clk);
#1;data_in = testData5[3978];
@(posedge clk);
#1;data_in = testData5[3979];
@(posedge clk);
#1;data_in = testData5[3980];
@(posedge clk);
#1;data_in = testData5[3981];
@(posedge clk);
#1;data_in = testData5[3982];
@(posedge clk);
#1;data_in = testData5[3983];
@(posedge clk);
#1;data_in = testData5[3984];
@(posedge clk);
#1;data_in = testData5[3985];
@(posedge clk);
#1;data_in = testData5[3986];
@(posedge clk);
#1;data_in = testData5[3987];
@(posedge clk);
#1;data_in = testData5[3988];
@(posedge clk);
#1;data_in = testData5[3989];
@(posedge clk);
#1;data_in = testData5[3990];
@(posedge clk);
#1;data_in = testData5[3991];
@(posedge clk);
#1;data_in = testData5[3992];
@(posedge clk);
#1;data_in = testData5[3993];
@(posedge clk);
#1;data_in = testData5[3994];
@(posedge clk);
#1;data_in = testData5[3995];
@(posedge clk);
#1;data_in = testData5[3996];
@(posedge clk);
#1;data_in = testData5[3997];
@(posedge clk);
#1;data_in = testData5[3998];
@(posedge clk);
#1;data_in = testData5[3999];
@(posedge clk);
#1;data_in = testData5[4000];
@(posedge clk);
#1;data_in = testData5[4001];
@(posedge clk);
#1;data_in = testData5[4002];
@(posedge clk);
#1;data_in = testData5[4003];
@(posedge clk);
#1;data_in = testData5[4004];
@(posedge clk);
#1;data_in = testData5[4005];
@(posedge clk);
#1;data_in = testData5[4006];
@(posedge clk);
#1;data_in = testData5[4007];
@(posedge clk);
#1;data_in = testData5[4008];
@(posedge clk);
#1;data_in = testData5[4009];
@(posedge clk);
#1;data_in = testData5[4010];
@(posedge clk);
#1;data_in = testData5[4011];
@(posedge clk);
#1;data_in = testData5[4012];
@(posedge clk);
#1;data_in = testData5[4013];
@(posedge clk);
#1;data_in = testData5[4014];
@(posedge clk);
#1;data_in = testData5[4015];
@(posedge clk);
#1;data_in = testData5[4016];
@(posedge clk);
#1;data_in = testData5[4017];
@(posedge clk);
#1;data_in = testData5[4018];
@(posedge clk);
#1;data_in = testData5[4019];
@(posedge clk);
#1;data_in = testData5[4020];
@(posedge clk);
#1;data_in = testData5[4021];
@(posedge clk);
#1;data_in = testData5[4022];
@(posedge clk);
#1;data_in = testData5[4023];
@(posedge clk);
#1;data_in = testData5[4024];
@(posedge clk);
#1;data_in = testData5[4025];
@(posedge clk);
#1;data_in = testData5[4026];
@(posedge clk);
#1;data_in = testData5[4027];
@(posedge clk);
#1;data_in = testData5[4028];
@(posedge clk);
#1;data_in = testData5[4029];
@(posedge clk);
#1;data_in = testData5[4030];
@(posedge clk);
#1;data_in = testData5[4031];
@(posedge clk);
#1;data_in = testData5[4032];
@(posedge clk);
#1;data_in = testData5[4033];
@(posedge clk);
#1;data_in = testData5[4034];
@(posedge clk);
#1;data_in = testData5[4035];
@(posedge clk);
#1;data_in = testData5[4036];
@(posedge clk);
#1;data_in = testData5[4037];
@(posedge clk);
#1;data_in = testData5[4038];
@(posedge clk);
#1;data_in = testData5[4039];
@(posedge clk);
#1;data_in = testData5[4040];
@(posedge clk);
#1;data_in = testData5[4041];
@(posedge clk);
#1;data_in = testData5[4042];
@(posedge clk);
#1;data_in = testData5[4043];
@(posedge clk);
#1;data_in = testData5[4044];
@(posedge clk);
#1;data_in = testData5[4045];
@(posedge clk);
#1;data_in = testData5[4046];
@(posedge clk);
#1;data_in = testData5[4047];
@(posedge clk);
#1;data_in = testData5[4048];
@(posedge clk);
#1;data_in = testData5[4049];
@(posedge clk);
#1;data_in = testData5[4050];
@(posedge clk);
#1;data_in = testData5[4051];
@(posedge clk);
#1;data_in = testData5[4052];
@(posedge clk);
#1;data_in = testData5[4053];
@(posedge clk);
#1;data_in = testData5[4054];
@(posedge clk);
#1;data_in = testData5[4055];
@(posedge clk);
#1;data_in = testData5[4056];
@(posedge clk);
#1;data_in = testData5[4057];
@(posedge clk);
#1;data_in = testData5[4058];
@(posedge clk);
#1;data_in = testData5[4059];
@(posedge clk);
#1;data_in = testData5[4060];
@(posedge clk);
#1;data_in = testData5[4061];
@(posedge clk);
#1;data_in = testData5[4062];
@(posedge clk);
#1;data_in = testData5[4063];
@(posedge clk);
#1;data_in = testData5[4064];
@(posedge clk);
#1;data_in = testData5[4065];
@(posedge clk);
#1;data_in = testData5[4066];
@(posedge clk);
#1;data_in = testData5[4067];
@(posedge clk);
#1;data_in = testData5[4068];
@(posedge clk);
#1;data_in = testData5[4069];
@(posedge clk);
#1;data_in = testData5[4070];
@(posedge clk);
#1;data_in = testData5[4071];
@(posedge clk);
#1;data_in = testData5[4072];
@(posedge clk);
#1;data_in = testData5[4073];
@(posedge clk);
#1;data_in = testData5[4074];
@(posedge clk);
#1;data_in = testData5[4075];
@(posedge clk);
#1;data_in = testData5[4076];
@(posedge clk);
#1;data_in = testData5[4077];
@(posedge clk);
#1;data_in = testData5[4078];
@(posedge clk);
#1;data_in = testData5[4079];
@(posedge clk);
#1;data_in = testData5[4080];
@(posedge clk);
#1;data_in = testData5[4081];
@(posedge clk);
#1;data_in = testData5[4082];
@(posedge clk);
#1;data_in = testData5[4083];
@(posedge clk);
#1;data_in = testData5[4084];
@(posedge clk);
#1;data_in = testData5[4085];
@(posedge clk);
#1;data_in = testData5[4086];
@(posedge clk);
#1;data_in = testData5[4087];
@(posedge clk);
#1;data_in = testData5[4088];
@(posedge clk);
#1;data_in = testData5[4089];
@(posedge clk);
#1;data_in = testData5[4090];
@(posedge clk);
#1;data_in = testData5[4091];
@(posedge clk);
#1;data_in = testData5[4092];
@(posedge clk);
#1;data_in = testData5[4093];
@(posedge clk);
#1;data_in = testData5[4094];
@(posedge clk);
#1;data_in = testData5[4095];
@(posedge clk);
#1;data_in = testData5[4096];
@(posedge clk);
#1;data_in = testData5[4097];
@(posedge clk);
#1;data_in = testData5[4098];
@(posedge clk);
#1;data_in = testData5[4099];
@(posedge clk);
#1;data_in = testData5[4100];
@(posedge clk);
#1;data_in = testData5[4101];
@(posedge clk);
#1;data_in = testData5[4102];
@(posedge clk);
#1;data_in = testData5[4103];
@(posedge clk);
#1;data_in = testData5[4104];
@(posedge clk);
#1;data_in = testData5[4105];
@(posedge clk);
#1;data_in = testData5[4106];
@(posedge clk);
#1;data_in = testData5[4107];
@(posedge clk);
#1;data_in = testData5[4108];
@(posedge clk);
#1;data_in = testData5[4109];
@(posedge clk);
#1;data_in = testData5[4110];
@(posedge clk);
#1;data_in = testData5[4111];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[4112]; 
@(posedge clk);
#1;data_in = testData5[4113];
@(posedge clk);
#1;data_in = testData5[4114];
@(posedge clk);
#1;data_in = testData5[4115];
@(posedge clk);
#1;data_in = testData5[4116];
@(posedge clk);
#1;data_in = testData5[4117];
@(posedge clk);
#1;data_in = testData5[4118];
@(posedge clk);
#1;data_in = testData5[4119];
@(posedge clk);
#1;data_in = testData5[4120];
@(posedge clk);
#1;data_in = testData5[4121];
@(posedge clk);
#1;data_in = testData5[4122];
@(posedge clk);
#1;data_in = testData5[4123];
@(posedge clk);
#1;data_in = testData5[4124];
@(posedge clk);
#1;data_in = testData5[4125];
@(posedge clk);
#1;data_in = testData5[4126];
@(posedge clk);
#1;data_in = testData5[4127];
@(posedge clk);
#1;data_in = testData5[4128];
@(posedge clk);
#1;data_in = testData5[4129];
@(posedge clk);
#1;data_in = testData5[4130];
@(posedge clk);
#1;data_in = testData5[4131];
@(posedge clk);
#1;data_in = testData5[4132];
@(posedge clk);
#1;data_in = testData5[4133];
@(posedge clk);
#1;data_in = testData5[4134];
@(posedge clk);
#1;data_in = testData5[4135];
@(posedge clk);
#1;data_in = testData5[4136];
@(posedge clk);
#1;data_in = testData5[4137];
@(posedge clk);
#1;data_in = testData5[4138];
@(posedge clk);
#1;data_in = testData5[4139];
@(posedge clk);
#1;data_in = testData5[4140];
@(posedge clk);
#1;data_in = testData5[4141];
@(posedge clk);
#1;data_in = testData5[4142];
@(posedge clk);
#1;data_in = testData5[4143];
@(posedge clk);
#1;data_in = testData5[4144];
@(posedge clk);
#1;data_in = testData5[4145];
@(posedge clk);
#1;data_in = testData5[4146];
@(posedge clk);
#1;data_in = testData5[4147];
@(posedge clk);
#1;data_in = testData5[4148];
@(posedge clk);
#1;data_in = testData5[4149];
@(posedge clk);
#1;data_in = testData5[4150];
@(posedge clk);
#1;data_in = testData5[4151];
@(posedge clk);
#1;data_in = testData5[4152];
@(posedge clk);
#1;data_in = testData5[4153];
@(posedge clk);
#1;data_in = testData5[4154];
@(posedge clk);
#1;data_in = testData5[4155];
@(posedge clk);
#1;data_in = testData5[4156];
@(posedge clk);
#1;data_in = testData5[4157];
@(posedge clk);
#1;data_in = testData5[4158];
@(posedge clk);
#1;data_in = testData5[4159];
@(posedge clk);
#1;data_in = testData5[4160];
@(posedge clk);
#1;data_in = testData5[4161];
@(posedge clk);
#1;data_in = testData5[4162];
@(posedge clk);
#1;data_in = testData5[4163];
@(posedge clk);
#1;data_in = testData5[4164];
@(posedge clk);
#1;data_in = testData5[4165];
@(posedge clk);
#1;data_in = testData5[4166];
@(posedge clk);
#1;data_in = testData5[4167];
@(posedge clk);
#1;data_in = testData5[4168];
@(posedge clk);
#1;data_in = testData5[4169];
@(posedge clk);
#1;data_in = testData5[4170];
@(posedge clk);
#1;data_in = testData5[4171];
@(posedge clk);
#1;data_in = testData5[4172];
@(posedge clk);
#1;data_in = testData5[4173];
@(posedge clk);
#1;data_in = testData5[4174];
@(posedge clk);
#1;data_in = testData5[4175];
@(posedge clk);
#1;data_in = testData5[4176];
@(posedge clk);
#1;data_in = testData5[4177];
@(posedge clk);
#1;data_in = testData5[4178];
@(posedge clk);
#1;data_in = testData5[4179];
@(posedge clk);
#1;data_in = testData5[4180];
@(posedge clk);
#1;data_in = testData5[4181];
@(posedge clk);
#1;data_in = testData5[4182];
@(posedge clk);
#1;data_in = testData5[4183];
@(posedge clk);
#1;data_in = testData5[4184];
@(posedge clk);
#1;data_in = testData5[4185];
@(posedge clk);
#1;data_in = testData5[4186];
@(posedge clk);
#1;data_in = testData5[4187];
@(posedge clk);
#1;data_in = testData5[4188];
@(posedge clk);
#1;data_in = testData5[4189];
@(posedge clk);
#1;data_in = testData5[4190];
@(posedge clk);
#1;data_in = testData5[4191];
@(posedge clk);
#1;data_in = testData5[4192];
@(posedge clk);
#1;data_in = testData5[4193];
@(posedge clk);
#1;data_in = testData5[4194];
@(posedge clk);
#1;data_in = testData5[4195];
@(posedge clk);
#1;data_in = testData5[4196];
@(posedge clk);
#1;data_in = testData5[4197];
@(posedge clk);
#1;data_in = testData5[4198];
@(posedge clk);
#1;data_in = testData5[4199];
@(posedge clk);
#1;data_in = testData5[4200];
@(posedge clk);
#1;data_in = testData5[4201];
@(posedge clk);
#1;data_in = testData5[4202];
@(posedge clk);
#1;data_in = testData5[4203];
@(posedge clk);
#1;data_in = testData5[4204];
@(posedge clk);
#1;data_in = testData5[4205];
@(posedge clk);
#1;data_in = testData5[4206];
@(posedge clk);
#1;data_in = testData5[4207];
@(posedge clk);
#1;data_in = testData5[4208];
@(posedge clk);
#1;data_in = testData5[4209];
@(posedge clk);
#1;data_in = testData5[4210];
@(posedge clk);
#1;data_in = testData5[4211];
@(posedge clk);
#1;data_in = testData5[4212];
@(posedge clk);
#1;data_in = testData5[4213];
@(posedge clk);
#1;data_in = testData5[4214];
@(posedge clk);
#1;data_in = testData5[4215];
@(posedge clk);
#1;data_in = testData5[4216];
@(posedge clk);
#1;data_in = testData5[4217];
@(posedge clk);
#1;data_in = testData5[4218];
@(posedge clk);
#1;data_in = testData5[4219];
@(posedge clk);
#1;data_in = testData5[4220];
@(posedge clk);
#1;data_in = testData5[4221];
@(posedge clk);
#1;data_in = testData5[4222];
@(posedge clk);
#1;data_in = testData5[4223];
@(posedge clk);
#1;data_in = testData5[4224];
@(posedge clk);
#1;data_in = testData5[4225];
@(posedge clk);
#1;data_in = testData5[4226];
@(posedge clk);
#1;data_in = testData5[4227];
@(posedge clk);
#1;data_in = testData5[4228];
@(posedge clk);
#1;data_in = testData5[4229];
@(posedge clk);
#1;data_in = testData5[4230];
@(posedge clk);
#1;data_in = testData5[4231];
@(posedge clk);
#1;data_in = testData5[4232];
@(posedge clk);
#1;data_in = testData5[4233];
@(posedge clk);
#1;data_in = testData5[4234];
@(posedge clk);
#1;data_in = testData5[4235];
@(posedge clk);
#1;data_in = testData5[4236];
@(posedge clk);
#1;data_in = testData5[4237];
@(posedge clk);
#1;data_in = testData5[4238];
@(posedge clk);
#1;data_in = testData5[4239];
@(posedge clk);
#1;data_in = testData5[4240];
@(posedge clk);
#1;data_in = testData5[4241];
@(posedge clk);
#1;data_in = testData5[4242];
@(posedge clk);
#1;data_in = testData5[4243];
@(posedge clk);
#1;data_in = testData5[4244];
@(posedge clk);
#1;data_in = testData5[4245];
@(posedge clk);
#1;data_in = testData5[4246];
@(posedge clk);
#1;data_in = testData5[4247];
@(posedge clk);
#1;data_in = testData5[4248];
@(posedge clk);
#1;data_in = testData5[4249];
@(posedge clk);
#1;data_in = testData5[4250];
@(posedge clk);
#1;data_in = testData5[4251];
@(posedge clk);
#1;data_in = testData5[4252];
@(posedge clk);
#1;data_in = testData5[4253];
@(posedge clk);
#1;data_in = testData5[4254];
@(posedge clk);
#1;data_in = testData5[4255];
@(posedge clk);
#1;data_in = testData5[4256];
@(posedge clk);
#1;data_in = testData5[4257];
@(posedge clk);
#1;data_in = testData5[4258];
@(posedge clk);
#1;data_in = testData5[4259];
@(posedge clk);
#1;data_in = testData5[4260];
@(posedge clk);
#1;data_in = testData5[4261];
@(posedge clk);
#1;data_in = testData5[4262];
@(posedge clk);
#1;data_in = testData5[4263];
@(posedge clk);
#1;data_in = testData5[4264];
@(posedge clk);
#1;data_in = testData5[4265];
@(posedge clk);
#1;data_in = testData5[4266];
@(posedge clk);
#1;data_in = testData5[4267];
@(posedge clk);
#1;data_in = testData5[4268];
@(posedge clk);
#1;data_in = testData5[4269];
@(posedge clk);
#1;data_in = testData5[4270];
@(posedge clk);
#1;data_in = testData5[4271];
@(posedge clk);
#1;data_in = testData5[4272];
@(posedge clk);
#1;data_in = testData5[4273];
@(posedge clk);
#1;data_in = testData5[4274];
@(posedge clk);
#1;data_in = testData5[4275];
@(posedge clk);
#1;data_in = testData5[4276];
@(posedge clk);
#1;data_in = testData5[4277];
@(posedge clk);
#1;data_in = testData5[4278];
@(posedge clk);
#1;data_in = testData5[4279];
@(posedge clk);
#1;data_in = testData5[4280];
@(posedge clk);
#1;data_in = testData5[4281];
@(posedge clk);
#1;data_in = testData5[4282];
@(posedge clk);
#1;data_in = testData5[4283];
@(posedge clk);
#1;data_in = testData5[4284];
@(posedge clk);
#1;data_in = testData5[4285];
@(posedge clk);
#1;data_in = testData5[4286];
@(posedge clk);
#1;data_in = testData5[4287];
@(posedge clk);
#1;data_in = testData5[4288];
@(posedge clk);
#1;data_in = testData5[4289];
@(posedge clk);
#1;data_in = testData5[4290];
@(posedge clk);
#1;data_in = testData5[4291];
@(posedge clk);
#1;data_in = testData5[4292];
@(posedge clk);
#1;data_in = testData5[4293];
@(posedge clk);
#1;data_in = testData5[4294];
@(posedge clk);
#1;data_in = testData5[4295];
@(posedge clk);
#1;data_in = testData5[4296];
@(posedge clk);
#1;data_in = testData5[4297];
@(posedge clk);
#1;data_in = testData5[4298];
@(posedge clk);
#1;data_in = testData5[4299];
@(posedge clk);
#1;data_in = testData5[4300];
@(posedge clk);
#1;data_in = testData5[4301];
@(posedge clk);
#1;data_in = testData5[4302];
@(posedge clk);
#1;data_in = testData5[4303];
@(posedge clk);
#1;data_in = testData5[4304];
@(posedge clk);
#1;data_in = testData5[4305];
@(posedge clk);
#1;data_in = testData5[4306];
@(posedge clk);
#1;data_in = testData5[4307];
@(posedge clk);
#1;data_in = testData5[4308];
@(posedge clk);
#1;data_in = testData5[4309];
@(posedge clk);
#1;data_in = testData5[4310];
@(posedge clk);
#1;data_in = testData5[4311];
@(posedge clk);
#1;data_in = testData5[4312];
@(posedge clk);
#1;data_in = testData5[4313];
@(posedge clk);
#1;data_in = testData5[4314];
@(posedge clk);
#1;data_in = testData5[4315];
@(posedge clk);
#1;data_in = testData5[4316];
@(posedge clk);
#1;data_in = testData5[4317];
@(posedge clk);
#1;data_in = testData5[4318];
@(posedge clk);
#1;data_in = testData5[4319];
@(posedge clk);
#1;data_in = testData5[4320];
@(posedge clk);
#1;data_in = testData5[4321];
@(posedge clk);
#1;data_in = testData5[4322];
@(posedge clk);
#1;data_in = testData5[4323];
@(posedge clk);
#1;data_in = testData5[4324];
@(posedge clk);
#1;data_in = testData5[4325];
@(posedge clk);
#1;data_in = testData5[4326];
@(posedge clk);
#1;data_in = testData5[4327];
@(posedge clk);
#1;data_in = testData5[4328];
@(posedge clk);
#1;data_in = testData5[4329];
@(posedge clk);
#1;data_in = testData5[4330];
@(posedge clk);
#1;data_in = testData5[4331];
@(posedge clk);
#1;data_in = testData5[4332];
@(posedge clk);
#1;data_in = testData5[4333];
@(posedge clk);
#1;data_in = testData5[4334];
@(posedge clk);
#1;data_in = testData5[4335];
@(posedge clk);
#1;data_in = testData5[4336];
@(posedge clk);
#1;data_in = testData5[4337];
@(posedge clk);
#1;data_in = testData5[4338];
@(posedge clk);
#1;data_in = testData5[4339];
@(posedge clk);
#1;data_in = testData5[4340];
@(posedge clk);
#1;data_in = testData5[4341];
@(posedge clk);
#1;data_in = testData5[4342];
@(posedge clk);
#1;data_in = testData5[4343];
@(posedge clk);
#1;data_in = testData5[4344];
@(posedge clk);
#1;data_in = testData5[4345];
@(posedge clk);
#1;data_in = testData5[4346];
@(posedge clk);
#1;data_in = testData5[4347];
@(posedge clk);
#1;data_in = testData5[4348];
@(posedge clk);
#1;data_in = testData5[4349];
@(posedge clk);
#1;data_in = testData5[4350];
@(posedge clk);
#1;data_in = testData5[4351];
@(posedge clk);
#1;data_in = testData5[4352];
@(posedge clk);
#1;data_in = testData5[4353];
@(posedge clk);
#1;data_in = testData5[4354];
@(posedge clk);
#1;data_in = testData5[4355];
@(posedge clk);
#1;data_in = testData5[4356];
@(posedge clk);
#1;data_in = testData5[4357];
@(posedge clk);
#1;data_in = testData5[4358];
@(posedge clk);
#1;data_in = testData5[4359];
@(posedge clk);
#1;data_in = testData5[4360];
@(posedge clk);
#1;data_in = testData5[4361];
@(posedge clk);
#1;data_in = testData5[4362];
@(posedge clk);
#1;data_in = testData5[4363];
@(posedge clk);
#1;data_in = testData5[4364];
@(posedge clk);
#1;data_in = testData5[4365];
@(posedge clk);
#1;data_in = testData5[4366];
@(posedge clk);
#1;data_in = testData5[4367];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[4368]; 
@(posedge clk);
#1;data_in = testData5[4369];
@(posedge clk);
#1;data_in = testData5[4370];
@(posedge clk);
#1;data_in = testData5[4371];
@(posedge clk);
#1;data_in = testData5[4372];
@(posedge clk);
#1;data_in = testData5[4373];
@(posedge clk);
#1;data_in = testData5[4374];
@(posedge clk);
#1;data_in = testData5[4375];
@(posedge clk);
#1;data_in = testData5[4376];
@(posedge clk);
#1;data_in = testData5[4377];
@(posedge clk);
#1;data_in = testData5[4378];
@(posedge clk);
#1;data_in = testData5[4379];
@(posedge clk);
#1;data_in = testData5[4380];
@(posedge clk);
#1;data_in = testData5[4381];
@(posedge clk);
#1;data_in = testData5[4382];
@(posedge clk);
#1;data_in = testData5[4383];
@(posedge clk);
#1;data_in = testData5[4384];
@(posedge clk);
#1;data_in = testData5[4385];
@(posedge clk);
#1;data_in = testData5[4386];
@(posedge clk);
#1;data_in = testData5[4387];
@(posedge clk);
#1;data_in = testData5[4388];
@(posedge clk);
#1;data_in = testData5[4389];
@(posedge clk);
#1;data_in = testData5[4390];
@(posedge clk);
#1;data_in = testData5[4391];
@(posedge clk);
#1;data_in = testData5[4392];
@(posedge clk);
#1;data_in = testData5[4393];
@(posedge clk);
#1;data_in = testData5[4394];
@(posedge clk);
#1;data_in = testData5[4395];
@(posedge clk);
#1;data_in = testData5[4396];
@(posedge clk);
#1;data_in = testData5[4397];
@(posedge clk);
#1;data_in = testData5[4398];
@(posedge clk);
#1;data_in = testData5[4399];
@(posedge clk);
#1;data_in = testData5[4400];
@(posedge clk);
#1;data_in = testData5[4401];
@(posedge clk);
#1;data_in = testData5[4402];
@(posedge clk);
#1;data_in = testData5[4403];
@(posedge clk);
#1;data_in = testData5[4404];
@(posedge clk);
#1;data_in = testData5[4405];
@(posedge clk);
#1;data_in = testData5[4406];
@(posedge clk);
#1;data_in = testData5[4407];
@(posedge clk);
#1;data_in = testData5[4408];
@(posedge clk);
#1;data_in = testData5[4409];
@(posedge clk);
#1;data_in = testData5[4410];
@(posedge clk);
#1;data_in = testData5[4411];
@(posedge clk);
#1;data_in = testData5[4412];
@(posedge clk);
#1;data_in = testData5[4413];
@(posedge clk);
#1;data_in = testData5[4414];
@(posedge clk);
#1;data_in = testData5[4415];
@(posedge clk);
#1;data_in = testData5[4416];
@(posedge clk);
#1;data_in = testData5[4417];
@(posedge clk);
#1;data_in = testData5[4418];
@(posedge clk);
#1;data_in = testData5[4419];
@(posedge clk);
#1;data_in = testData5[4420];
@(posedge clk);
#1;data_in = testData5[4421];
@(posedge clk);
#1;data_in = testData5[4422];
@(posedge clk);
#1;data_in = testData5[4423];
@(posedge clk);
#1;data_in = testData5[4424];
@(posedge clk);
#1;data_in = testData5[4425];
@(posedge clk);
#1;data_in = testData5[4426];
@(posedge clk);
#1;data_in = testData5[4427];
@(posedge clk);
#1;data_in = testData5[4428];
@(posedge clk);
#1;data_in = testData5[4429];
@(posedge clk);
#1;data_in = testData5[4430];
@(posedge clk);
#1;data_in = testData5[4431];
@(posedge clk);
#1;data_in = testData5[4432];
@(posedge clk);
#1;data_in = testData5[4433];
@(posedge clk);
#1;data_in = testData5[4434];
@(posedge clk);
#1;data_in = testData5[4435];
@(posedge clk);
#1;data_in = testData5[4436];
@(posedge clk);
#1;data_in = testData5[4437];
@(posedge clk);
#1;data_in = testData5[4438];
@(posedge clk);
#1;data_in = testData5[4439];
@(posedge clk);
#1;data_in = testData5[4440];
@(posedge clk);
#1;data_in = testData5[4441];
@(posedge clk);
#1;data_in = testData5[4442];
@(posedge clk);
#1;data_in = testData5[4443];
@(posedge clk);
#1;data_in = testData5[4444];
@(posedge clk);
#1;data_in = testData5[4445];
@(posedge clk);
#1;data_in = testData5[4446];
@(posedge clk);
#1;data_in = testData5[4447];
@(posedge clk);
#1;data_in = testData5[4448];
@(posedge clk);
#1;data_in = testData5[4449];
@(posedge clk);
#1;data_in = testData5[4450];
@(posedge clk);
#1;data_in = testData5[4451];
@(posedge clk);
#1;data_in = testData5[4452];
@(posedge clk);
#1;data_in = testData5[4453];
@(posedge clk);
#1;data_in = testData5[4454];
@(posedge clk);
#1;data_in = testData5[4455];
@(posedge clk);
#1;data_in = testData5[4456];
@(posedge clk);
#1;data_in = testData5[4457];
@(posedge clk);
#1;data_in = testData5[4458];
@(posedge clk);
#1;data_in = testData5[4459];
@(posedge clk);
#1;data_in = testData5[4460];
@(posedge clk);
#1;data_in = testData5[4461];
@(posedge clk);
#1;data_in = testData5[4462];
@(posedge clk);
#1;data_in = testData5[4463];
@(posedge clk);
#1;data_in = testData5[4464];
@(posedge clk);
#1;data_in = testData5[4465];
@(posedge clk);
#1;data_in = testData5[4466];
@(posedge clk);
#1;data_in = testData5[4467];
@(posedge clk);
#1;data_in = testData5[4468];
@(posedge clk);
#1;data_in = testData5[4469];
@(posedge clk);
#1;data_in = testData5[4470];
@(posedge clk);
#1;data_in = testData5[4471];
@(posedge clk);
#1;data_in = testData5[4472];
@(posedge clk);
#1;data_in = testData5[4473];
@(posedge clk);
#1;data_in = testData5[4474];
@(posedge clk);
#1;data_in = testData5[4475];
@(posedge clk);
#1;data_in = testData5[4476];
@(posedge clk);
#1;data_in = testData5[4477];
@(posedge clk);
#1;data_in = testData5[4478];
@(posedge clk);
#1;data_in = testData5[4479];
@(posedge clk);
#1;data_in = testData5[4480];
@(posedge clk);
#1;data_in = testData5[4481];
@(posedge clk);
#1;data_in = testData5[4482];
@(posedge clk);
#1;data_in = testData5[4483];
@(posedge clk);
#1;data_in = testData5[4484];
@(posedge clk);
#1;data_in = testData5[4485];
@(posedge clk);
#1;data_in = testData5[4486];
@(posedge clk);
#1;data_in = testData5[4487];
@(posedge clk);
#1;data_in = testData5[4488];
@(posedge clk);
#1;data_in = testData5[4489];
@(posedge clk);
#1;data_in = testData5[4490];
@(posedge clk);
#1;data_in = testData5[4491];
@(posedge clk);
#1;data_in = testData5[4492];
@(posedge clk);
#1;data_in = testData5[4493];
@(posedge clk);
#1;data_in = testData5[4494];
@(posedge clk);
#1;data_in = testData5[4495];
@(posedge clk);
#1;data_in = testData5[4496];
@(posedge clk);
#1;data_in = testData5[4497];
@(posedge clk);
#1;data_in = testData5[4498];
@(posedge clk);
#1;data_in = testData5[4499];
@(posedge clk);
#1;data_in = testData5[4500];
@(posedge clk);
#1;data_in = testData5[4501];
@(posedge clk);
#1;data_in = testData5[4502];
@(posedge clk);
#1;data_in = testData5[4503];
@(posedge clk);
#1;data_in = testData5[4504];
@(posedge clk);
#1;data_in = testData5[4505];
@(posedge clk);
#1;data_in = testData5[4506];
@(posedge clk);
#1;data_in = testData5[4507];
@(posedge clk);
#1;data_in = testData5[4508];
@(posedge clk);
#1;data_in = testData5[4509];
@(posedge clk);
#1;data_in = testData5[4510];
@(posedge clk);
#1;data_in = testData5[4511];
@(posedge clk);
#1;data_in = testData5[4512];
@(posedge clk);
#1;data_in = testData5[4513];
@(posedge clk);
#1;data_in = testData5[4514];
@(posedge clk);
#1;data_in = testData5[4515];
@(posedge clk);
#1;data_in = testData5[4516];
@(posedge clk);
#1;data_in = testData5[4517];
@(posedge clk);
#1;data_in = testData5[4518];
@(posedge clk);
#1;data_in = testData5[4519];
@(posedge clk);
#1;data_in = testData5[4520];
@(posedge clk);
#1;data_in = testData5[4521];
@(posedge clk);
#1;data_in = testData5[4522];
@(posedge clk);
#1;data_in = testData5[4523];
@(posedge clk);
#1;data_in = testData5[4524];
@(posedge clk);
#1;data_in = testData5[4525];
@(posedge clk);
#1;data_in = testData5[4526];
@(posedge clk);
#1;data_in = testData5[4527];
@(posedge clk);
#1;data_in = testData5[4528];
@(posedge clk);
#1;data_in = testData5[4529];
@(posedge clk);
#1;data_in = testData5[4530];
@(posedge clk);
#1;data_in = testData5[4531];
@(posedge clk);
#1;data_in = testData5[4532];
@(posedge clk);
#1;data_in = testData5[4533];
@(posedge clk);
#1;data_in = testData5[4534];
@(posedge clk);
#1;data_in = testData5[4535];
@(posedge clk);
#1;data_in = testData5[4536];
@(posedge clk);
#1;data_in = testData5[4537];
@(posedge clk);
#1;data_in = testData5[4538];
@(posedge clk);
#1;data_in = testData5[4539];
@(posedge clk);
#1;data_in = testData5[4540];
@(posedge clk);
#1;data_in = testData5[4541];
@(posedge clk);
#1;data_in = testData5[4542];
@(posedge clk);
#1;data_in = testData5[4543];
@(posedge clk);
#1;data_in = testData5[4544];
@(posedge clk);
#1;data_in = testData5[4545];
@(posedge clk);
#1;data_in = testData5[4546];
@(posedge clk);
#1;data_in = testData5[4547];
@(posedge clk);
#1;data_in = testData5[4548];
@(posedge clk);
#1;data_in = testData5[4549];
@(posedge clk);
#1;data_in = testData5[4550];
@(posedge clk);
#1;data_in = testData5[4551];
@(posedge clk);
#1;data_in = testData5[4552];
@(posedge clk);
#1;data_in = testData5[4553];
@(posedge clk);
#1;data_in = testData5[4554];
@(posedge clk);
#1;data_in = testData5[4555];
@(posedge clk);
#1;data_in = testData5[4556];
@(posedge clk);
#1;data_in = testData5[4557];
@(posedge clk);
#1;data_in = testData5[4558];
@(posedge clk);
#1;data_in = testData5[4559];
@(posedge clk);
#1;data_in = testData5[4560];
@(posedge clk);
#1;data_in = testData5[4561];
@(posedge clk);
#1;data_in = testData5[4562];
@(posedge clk);
#1;data_in = testData5[4563];
@(posedge clk);
#1;data_in = testData5[4564];
@(posedge clk);
#1;data_in = testData5[4565];
@(posedge clk);
#1;data_in = testData5[4566];
@(posedge clk);
#1;data_in = testData5[4567];
@(posedge clk);
#1;data_in = testData5[4568];
@(posedge clk);
#1;data_in = testData5[4569];
@(posedge clk);
#1;data_in = testData5[4570];
@(posedge clk);
#1;data_in = testData5[4571];
@(posedge clk);
#1;data_in = testData5[4572];
@(posedge clk);
#1;data_in = testData5[4573];
@(posedge clk);
#1;data_in = testData5[4574];
@(posedge clk);
#1;data_in = testData5[4575];
@(posedge clk);
#1;data_in = testData5[4576];
@(posedge clk);
#1;data_in = testData5[4577];
@(posedge clk);
#1;data_in = testData5[4578];
@(posedge clk);
#1;data_in = testData5[4579];
@(posedge clk);
#1;data_in = testData5[4580];
@(posedge clk);
#1;data_in = testData5[4581];
@(posedge clk);
#1;data_in = testData5[4582];
@(posedge clk);
#1;data_in = testData5[4583];
@(posedge clk);
#1;data_in = testData5[4584];
@(posedge clk);
#1;data_in = testData5[4585];
@(posedge clk);
#1;data_in = testData5[4586];
@(posedge clk);
#1;data_in = testData5[4587];
@(posedge clk);
#1;data_in = testData5[4588];
@(posedge clk);
#1;data_in = testData5[4589];
@(posedge clk);
#1;data_in = testData5[4590];
@(posedge clk);
#1;data_in = testData5[4591];
@(posedge clk);
#1;data_in = testData5[4592];
@(posedge clk);
#1;data_in = testData5[4593];
@(posedge clk);
#1;data_in = testData5[4594];
@(posedge clk);
#1;data_in = testData5[4595];
@(posedge clk);
#1;data_in = testData5[4596];
@(posedge clk);
#1;data_in = testData5[4597];
@(posedge clk);
#1;data_in = testData5[4598];
@(posedge clk);
#1;data_in = testData5[4599];
@(posedge clk);
#1;data_in = testData5[4600];
@(posedge clk);
#1;data_in = testData5[4601];
@(posedge clk);
#1;data_in = testData5[4602];
@(posedge clk);
#1;data_in = testData5[4603];
@(posedge clk);
#1;data_in = testData5[4604];
@(posedge clk);
#1;data_in = testData5[4605];
@(posedge clk);
#1;data_in = testData5[4606];
@(posedge clk);
#1;data_in = testData5[4607];
@(posedge clk);
#1;data_in = testData5[4608];
@(posedge clk);
#1;data_in = testData5[4609];
@(posedge clk);
#1;data_in = testData5[4610];
@(posedge clk);
#1;data_in = testData5[4611];
@(posedge clk);
#1;data_in = testData5[4612];
@(posedge clk);
#1;data_in = testData5[4613];
@(posedge clk);
#1;data_in = testData5[4614];
@(posedge clk);
#1;data_in = testData5[4615];
@(posedge clk);
#1;data_in = testData5[4616];
@(posedge clk);
#1;data_in = testData5[4617];
@(posedge clk);
#1;data_in = testData5[4618];
@(posedge clk);
#1;data_in = testData5[4619];
@(posedge clk);
#1;data_in = testData5[4620];
@(posedge clk);
#1;data_in = testData5[4621];
@(posedge clk);
#1;data_in = testData5[4622];
@(posedge clk);
#1;data_in = testData5[4623];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[4624]; 
@(posedge clk);
#1;data_in = testData5[4625];
@(posedge clk);
#1;data_in = testData5[4626];
@(posedge clk);
#1;data_in = testData5[4627];
@(posedge clk);
#1;data_in = testData5[4628];
@(posedge clk);
#1;data_in = testData5[4629];
@(posedge clk);
#1;data_in = testData5[4630];
@(posedge clk);
#1;data_in = testData5[4631];
@(posedge clk);
#1;data_in = testData5[4632];
@(posedge clk);
#1;data_in = testData5[4633];
@(posedge clk);
#1;data_in = testData5[4634];
@(posedge clk);
#1;data_in = testData5[4635];
@(posedge clk);
#1;data_in = testData5[4636];
@(posedge clk);
#1;data_in = testData5[4637];
@(posedge clk);
#1;data_in = testData5[4638];
@(posedge clk);
#1;data_in = testData5[4639];
@(posedge clk);
#1;data_in = testData5[4640];
@(posedge clk);
#1;data_in = testData5[4641];
@(posedge clk);
#1;data_in = testData5[4642];
@(posedge clk);
#1;data_in = testData5[4643];
@(posedge clk);
#1;data_in = testData5[4644];
@(posedge clk);
#1;data_in = testData5[4645];
@(posedge clk);
#1;data_in = testData5[4646];
@(posedge clk);
#1;data_in = testData5[4647];
@(posedge clk);
#1;data_in = testData5[4648];
@(posedge clk);
#1;data_in = testData5[4649];
@(posedge clk);
#1;data_in = testData5[4650];
@(posedge clk);
#1;data_in = testData5[4651];
@(posedge clk);
#1;data_in = testData5[4652];
@(posedge clk);
#1;data_in = testData5[4653];
@(posedge clk);
#1;data_in = testData5[4654];
@(posedge clk);
#1;data_in = testData5[4655];
@(posedge clk);
#1;data_in = testData5[4656];
@(posedge clk);
#1;data_in = testData5[4657];
@(posedge clk);
#1;data_in = testData5[4658];
@(posedge clk);
#1;data_in = testData5[4659];
@(posedge clk);
#1;data_in = testData5[4660];
@(posedge clk);
#1;data_in = testData5[4661];
@(posedge clk);
#1;data_in = testData5[4662];
@(posedge clk);
#1;data_in = testData5[4663];
@(posedge clk);
#1;data_in = testData5[4664];
@(posedge clk);
#1;data_in = testData5[4665];
@(posedge clk);
#1;data_in = testData5[4666];
@(posedge clk);
#1;data_in = testData5[4667];
@(posedge clk);
#1;data_in = testData5[4668];
@(posedge clk);
#1;data_in = testData5[4669];
@(posedge clk);
#1;data_in = testData5[4670];
@(posedge clk);
#1;data_in = testData5[4671];
@(posedge clk);
#1;data_in = testData5[4672];
@(posedge clk);
#1;data_in = testData5[4673];
@(posedge clk);
#1;data_in = testData5[4674];
@(posedge clk);
#1;data_in = testData5[4675];
@(posedge clk);
#1;data_in = testData5[4676];
@(posedge clk);
#1;data_in = testData5[4677];
@(posedge clk);
#1;data_in = testData5[4678];
@(posedge clk);
#1;data_in = testData5[4679];
@(posedge clk);
#1;data_in = testData5[4680];
@(posedge clk);
#1;data_in = testData5[4681];
@(posedge clk);
#1;data_in = testData5[4682];
@(posedge clk);
#1;data_in = testData5[4683];
@(posedge clk);
#1;data_in = testData5[4684];
@(posedge clk);
#1;data_in = testData5[4685];
@(posedge clk);
#1;data_in = testData5[4686];
@(posedge clk);
#1;data_in = testData5[4687];
@(posedge clk);
#1;data_in = testData5[4688];
@(posedge clk);
#1;data_in = testData5[4689];
@(posedge clk);
#1;data_in = testData5[4690];
@(posedge clk);
#1;data_in = testData5[4691];
@(posedge clk);
#1;data_in = testData5[4692];
@(posedge clk);
#1;data_in = testData5[4693];
@(posedge clk);
#1;data_in = testData5[4694];
@(posedge clk);
#1;data_in = testData5[4695];
@(posedge clk);
#1;data_in = testData5[4696];
@(posedge clk);
#1;data_in = testData5[4697];
@(posedge clk);
#1;data_in = testData5[4698];
@(posedge clk);
#1;data_in = testData5[4699];
@(posedge clk);
#1;data_in = testData5[4700];
@(posedge clk);
#1;data_in = testData5[4701];
@(posedge clk);
#1;data_in = testData5[4702];
@(posedge clk);
#1;data_in = testData5[4703];
@(posedge clk);
#1;data_in = testData5[4704];
@(posedge clk);
#1;data_in = testData5[4705];
@(posedge clk);
#1;data_in = testData5[4706];
@(posedge clk);
#1;data_in = testData5[4707];
@(posedge clk);
#1;data_in = testData5[4708];
@(posedge clk);
#1;data_in = testData5[4709];
@(posedge clk);
#1;data_in = testData5[4710];
@(posedge clk);
#1;data_in = testData5[4711];
@(posedge clk);
#1;data_in = testData5[4712];
@(posedge clk);
#1;data_in = testData5[4713];
@(posedge clk);
#1;data_in = testData5[4714];
@(posedge clk);
#1;data_in = testData5[4715];
@(posedge clk);
#1;data_in = testData5[4716];
@(posedge clk);
#1;data_in = testData5[4717];
@(posedge clk);
#1;data_in = testData5[4718];
@(posedge clk);
#1;data_in = testData5[4719];
@(posedge clk);
#1;data_in = testData5[4720];
@(posedge clk);
#1;data_in = testData5[4721];
@(posedge clk);
#1;data_in = testData5[4722];
@(posedge clk);
#1;data_in = testData5[4723];
@(posedge clk);
#1;data_in = testData5[4724];
@(posedge clk);
#1;data_in = testData5[4725];
@(posedge clk);
#1;data_in = testData5[4726];
@(posedge clk);
#1;data_in = testData5[4727];
@(posedge clk);
#1;data_in = testData5[4728];
@(posedge clk);
#1;data_in = testData5[4729];
@(posedge clk);
#1;data_in = testData5[4730];
@(posedge clk);
#1;data_in = testData5[4731];
@(posedge clk);
#1;data_in = testData5[4732];
@(posedge clk);
#1;data_in = testData5[4733];
@(posedge clk);
#1;data_in = testData5[4734];
@(posedge clk);
#1;data_in = testData5[4735];
@(posedge clk);
#1;data_in = testData5[4736];
@(posedge clk);
#1;data_in = testData5[4737];
@(posedge clk);
#1;data_in = testData5[4738];
@(posedge clk);
#1;data_in = testData5[4739];
@(posedge clk);
#1;data_in = testData5[4740];
@(posedge clk);
#1;data_in = testData5[4741];
@(posedge clk);
#1;data_in = testData5[4742];
@(posedge clk);
#1;data_in = testData5[4743];
@(posedge clk);
#1;data_in = testData5[4744];
@(posedge clk);
#1;data_in = testData5[4745];
@(posedge clk);
#1;data_in = testData5[4746];
@(posedge clk);
#1;data_in = testData5[4747];
@(posedge clk);
#1;data_in = testData5[4748];
@(posedge clk);
#1;data_in = testData5[4749];
@(posedge clk);
#1;data_in = testData5[4750];
@(posedge clk);
#1;data_in = testData5[4751];
@(posedge clk);
#1;data_in = testData5[4752];
@(posedge clk);
#1;data_in = testData5[4753];
@(posedge clk);
#1;data_in = testData5[4754];
@(posedge clk);
#1;data_in = testData5[4755];
@(posedge clk);
#1;data_in = testData5[4756];
@(posedge clk);
#1;data_in = testData5[4757];
@(posedge clk);
#1;data_in = testData5[4758];
@(posedge clk);
#1;data_in = testData5[4759];
@(posedge clk);
#1;data_in = testData5[4760];
@(posedge clk);
#1;data_in = testData5[4761];
@(posedge clk);
#1;data_in = testData5[4762];
@(posedge clk);
#1;data_in = testData5[4763];
@(posedge clk);
#1;data_in = testData5[4764];
@(posedge clk);
#1;data_in = testData5[4765];
@(posedge clk);
#1;data_in = testData5[4766];
@(posedge clk);
#1;data_in = testData5[4767];
@(posedge clk);
#1;data_in = testData5[4768];
@(posedge clk);
#1;data_in = testData5[4769];
@(posedge clk);
#1;data_in = testData5[4770];
@(posedge clk);
#1;data_in = testData5[4771];
@(posedge clk);
#1;data_in = testData5[4772];
@(posedge clk);
#1;data_in = testData5[4773];
@(posedge clk);
#1;data_in = testData5[4774];
@(posedge clk);
#1;data_in = testData5[4775];
@(posedge clk);
#1;data_in = testData5[4776];
@(posedge clk);
#1;data_in = testData5[4777];
@(posedge clk);
#1;data_in = testData5[4778];
@(posedge clk);
#1;data_in = testData5[4779];
@(posedge clk);
#1;data_in = testData5[4780];
@(posedge clk);
#1;data_in = testData5[4781];
@(posedge clk);
#1;data_in = testData5[4782];
@(posedge clk);
#1;data_in = testData5[4783];
@(posedge clk);
#1;data_in = testData5[4784];
@(posedge clk);
#1;data_in = testData5[4785];
@(posedge clk);
#1;data_in = testData5[4786];
@(posedge clk);
#1;data_in = testData5[4787];
@(posedge clk);
#1;data_in = testData5[4788];
@(posedge clk);
#1;data_in = testData5[4789];
@(posedge clk);
#1;data_in = testData5[4790];
@(posedge clk);
#1;data_in = testData5[4791];
@(posedge clk);
#1;data_in = testData5[4792];
@(posedge clk);
#1;data_in = testData5[4793];
@(posedge clk);
#1;data_in = testData5[4794];
@(posedge clk);
#1;data_in = testData5[4795];
@(posedge clk);
#1;data_in = testData5[4796];
@(posedge clk);
#1;data_in = testData5[4797];
@(posedge clk);
#1;data_in = testData5[4798];
@(posedge clk);
#1;data_in = testData5[4799];
@(posedge clk);
#1;data_in = testData5[4800];
@(posedge clk);
#1;data_in = testData5[4801];
@(posedge clk);
#1;data_in = testData5[4802];
@(posedge clk);
#1;data_in = testData5[4803];
@(posedge clk);
#1;data_in = testData5[4804];
@(posedge clk);
#1;data_in = testData5[4805];
@(posedge clk);
#1;data_in = testData5[4806];
@(posedge clk);
#1;data_in = testData5[4807];
@(posedge clk);
#1;data_in = testData5[4808];
@(posedge clk);
#1;data_in = testData5[4809];
@(posedge clk);
#1;data_in = testData5[4810];
@(posedge clk);
#1;data_in = testData5[4811];
@(posedge clk);
#1;data_in = testData5[4812];
@(posedge clk);
#1;data_in = testData5[4813];
@(posedge clk);
#1;data_in = testData5[4814];
@(posedge clk);
#1;data_in = testData5[4815];
@(posedge clk);
#1;data_in = testData5[4816];
@(posedge clk);
#1;data_in = testData5[4817];
@(posedge clk);
#1;data_in = testData5[4818];
@(posedge clk);
#1;data_in = testData5[4819];
@(posedge clk);
#1;data_in = testData5[4820];
@(posedge clk);
#1;data_in = testData5[4821];
@(posedge clk);
#1;data_in = testData5[4822];
@(posedge clk);
#1;data_in = testData5[4823];
@(posedge clk);
#1;data_in = testData5[4824];
@(posedge clk);
#1;data_in = testData5[4825];
@(posedge clk);
#1;data_in = testData5[4826];
@(posedge clk);
#1;data_in = testData5[4827];
@(posedge clk);
#1;data_in = testData5[4828];
@(posedge clk);
#1;data_in = testData5[4829];
@(posedge clk);
#1;data_in = testData5[4830];
@(posedge clk);
#1;data_in = testData5[4831];
@(posedge clk);
#1;data_in = testData5[4832];
@(posedge clk);
#1;data_in = testData5[4833];
@(posedge clk);
#1;data_in = testData5[4834];
@(posedge clk);
#1;data_in = testData5[4835];
@(posedge clk);
#1;data_in = testData5[4836];
@(posedge clk);
#1;data_in = testData5[4837];
@(posedge clk);
#1;data_in = testData5[4838];
@(posedge clk);
#1;data_in = testData5[4839];
@(posedge clk);
#1;data_in = testData5[4840];
@(posedge clk);
#1;data_in = testData5[4841];
@(posedge clk);
#1;data_in = testData5[4842];
@(posedge clk);
#1;data_in = testData5[4843];
@(posedge clk);
#1;data_in = testData5[4844];
@(posedge clk);
#1;data_in = testData5[4845];
@(posedge clk);
#1;data_in = testData5[4846];
@(posedge clk);
#1;data_in = testData5[4847];
@(posedge clk);
#1;data_in = testData5[4848];
@(posedge clk);
#1;data_in = testData5[4849];
@(posedge clk);
#1;data_in = testData5[4850];
@(posedge clk);
#1;data_in = testData5[4851];
@(posedge clk);
#1;data_in = testData5[4852];
@(posedge clk);
#1;data_in = testData5[4853];
@(posedge clk);
#1;data_in = testData5[4854];
@(posedge clk);
#1;data_in = testData5[4855];
@(posedge clk);
#1;data_in = testData5[4856];
@(posedge clk);
#1;data_in = testData5[4857];
@(posedge clk);
#1;data_in = testData5[4858];
@(posedge clk);
#1;data_in = testData5[4859];
@(posedge clk);
#1;data_in = testData5[4860];
@(posedge clk);
#1;data_in = testData5[4861];
@(posedge clk);
#1;data_in = testData5[4862];
@(posedge clk);
#1;data_in = testData5[4863];
@(posedge clk);
#1;data_in = testData5[4864];
@(posedge clk);
#1;data_in = testData5[4865];
@(posedge clk);
#1;data_in = testData5[4866];
@(posedge clk);
#1;data_in = testData5[4867];
@(posedge clk);
#1;data_in = testData5[4868];
@(posedge clk);
#1;data_in = testData5[4869];
@(posedge clk);
#1;data_in = testData5[4870];
@(posedge clk);
#1;data_in = testData5[4871];
@(posedge clk);
#1;data_in = testData5[4872];
@(posedge clk);
#1;data_in = testData5[4873];
@(posedge clk);
#1;data_in = testData5[4874];
@(posedge clk);
#1;data_in = testData5[4875];
@(posedge clk);
#1;data_in = testData5[4876];
@(posedge clk);
#1;data_in = testData5[4877];
@(posedge clk);
#1;data_in = testData5[4878];
@(posedge clk);
#1;data_in = testData5[4879];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[4880]; 
@(posedge clk);
#1;data_in = testData5[4881];
@(posedge clk);
#1;data_in = testData5[4882];
@(posedge clk);
#1;data_in = testData5[4883];
@(posedge clk);
#1;data_in = testData5[4884];
@(posedge clk);
#1;data_in = testData5[4885];
@(posedge clk);
#1;data_in = testData5[4886];
@(posedge clk);
#1;data_in = testData5[4887];
@(posedge clk);
#1;data_in = testData5[4888];
@(posedge clk);
#1;data_in = testData5[4889];
@(posedge clk);
#1;data_in = testData5[4890];
@(posedge clk);
#1;data_in = testData5[4891];
@(posedge clk);
#1;data_in = testData5[4892];
@(posedge clk);
#1;data_in = testData5[4893];
@(posedge clk);
#1;data_in = testData5[4894];
@(posedge clk);
#1;data_in = testData5[4895];
@(posedge clk);
#1;data_in = testData5[4896];
@(posedge clk);
#1;data_in = testData5[4897];
@(posedge clk);
#1;data_in = testData5[4898];
@(posedge clk);
#1;data_in = testData5[4899];
@(posedge clk);
#1;data_in = testData5[4900];
@(posedge clk);
#1;data_in = testData5[4901];
@(posedge clk);
#1;data_in = testData5[4902];
@(posedge clk);
#1;data_in = testData5[4903];
@(posedge clk);
#1;data_in = testData5[4904];
@(posedge clk);
#1;data_in = testData5[4905];
@(posedge clk);
#1;data_in = testData5[4906];
@(posedge clk);
#1;data_in = testData5[4907];
@(posedge clk);
#1;data_in = testData5[4908];
@(posedge clk);
#1;data_in = testData5[4909];
@(posedge clk);
#1;data_in = testData5[4910];
@(posedge clk);
#1;data_in = testData5[4911];
@(posedge clk);
#1;data_in = testData5[4912];
@(posedge clk);
#1;data_in = testData5[4913];
@(posedge clk);
#1;data_in = testData5[4914];
@(posedge clk);
#1;data_in = testData5[4915];
@(posedge clk);
#1;data_in = testData5[4916];
@(posedge clk);
#1;data_in = testData5[4917];
@(posedge clk);
#1;data_in = testData5[4918];
@(posedge clk);
#1;data_in = testData5[4919];
@(posedge clk);
#1;data_in = testData5[4920];
@(posedge clk);
#1;data_in = testData5[4921];
@(posedge clk);
#1;data_in = testData5[4922];
@(posedge clk);
#1;data_in = testData5[4923];
@(posedge clk);
#1;data_in = testData5[4924];
@(posedge clk);
#1;data_in = testData5[4925];
@(posedge clk);
#1;data_in = testData5[4926];
@(posedge clk);
#1;data_in = testData5[4927];
@(posedge clk);
#1;data_in = testData5[4928];
@(posedge clk);
#1;data_in = testData5[4929];
@(posedge clk);
#1;data_in = testData5[4930];
@(posedge clk);
#1;data_in = testData5[4931];
@(posedge clk);
#1;data_in = testData5[4932];
@(posedge clk);
#1;data_in = testData5[4933];
@(posedge clk);
#1;data_in = testData5[4934];
@(posedge clk);
#1;data_in = testData5[4935];
@(posedge clk);
#1;data_in = testData5[4936];
@(posedge clk);
#1;data_in = testData5[4937];
@(posedge clk);
#1;data_in = testData5[4938];
@(posedge clk);
#1;data_in = testData5[4939];
@(posedge clk);
#1;data_in = testData5[4940];
@(posedge clk);
#1;data_in = testData5[4941];
@(posedge clk);
#1;data_in = testData5[4942];
@(posedge clk);
#1;data_in = testData5[4943];
@(posedge clk);
#1;data_in = testData5[4944];
@(posedge clk);
#1;data_in = testData5[4945];
@(posedge clk);
#1;data_in = testData5[4946];
@(posedge clk);
#1;data_in = testData5[4947];
@(posedge clk);
#1;data_in = testData5[4948];
@(posedge clk);
#1;data_in = testData5[4949];
@(posedge clk);
#1;data_in = testData5[4950];
@(posedge clk);
#1;data_in = testData5[4951];
@(posedge clk);
#1;data_in = testData5[4952];
@(posedge clk);
#1;data_in = testData5[4953];
@(posedge clk);
#1;data_in = testData5[4954];
@(posedge clk);
#1;data_in = testData5[4955];
@(posedge clk);
#1;data_in = testData5[4956];
@(posedge clk);
#1;data_in = testData5[4957];
@(posedge clk);
#1;data_in = testData5[4958];
@(posedge clk);
#1;data_in = testData5[4959];
@(posedge clk);
#1;data_in = testData5[4960];
@(posedge clk);
#1;data_in = testData5[4961];
@(posedge clk);
#1;data_in = testData5[4962];
@(posedge clk);
#1;data_in = testData5[4963];
@(posedge clk);
#1;data_in = testData5[4964];
@(posedge clk);
#1;data_in = testData5[4965];
@(posedge clk);
#1;data_in = testData5[4966];
@(posedge clk);
#1;data_in = testData5[4967];
@(posedge clk);
#1;data_in = testData5[4968];
@(posedge clk);
#1;data_in = testData5[4969];
@(posedge clk);
#1;data_in = testData5[4970];
@(posedge clk);
#1;data_in = testData5[4971];
@(posedge clk);
#1;data_in = testData5[4972];
@(posedge clk);
#1;data_in = testData5[4973];
@(posedge clk);
#1;data_in = testData5[4974];
@(posedge clk);
#1;data_in = testData5[4975];
@(posedge clk);
#1;data_in = testData5[4976];
@(posedge clk);
#1;data_in = testData5[4977];
@(posedge clk);
#1;data_in = testData5[4978];
@(posedge clk);
#1;data_in = testData5[4979];
@(posedge clk);
#1;data_in = testData5[4980];
@(posedge clk);
#1;data_in = testData5[4981];
@(posedge clk);
#1;data_in = testData5[4982];
@(posedge clk);
#1;data_in = testData5[4983];
@(posedge clk);
#1;data_in = testData5[4984];
@(posedge clk);
#1;data_in = testData5[4985];
@(posedge clk);
#1;data_in = testData5[4986];
@(posedge clk);
#1;data_in = testData5[4987];
@(posedge clk);
#1;data_in = testData5[4988];
@(posedge clk);
#1;data_in = testData5[4989];
@(posedge clk);
#1;data_in = testData5[4990];
@(posedge clk);
#1;data_in = testData5[4991];
@(posedge clk);
#1;data_in = testData5[4992];
@(posedge clk);
#1;data_in = testData5[4993];
@(posedge clk);
#1;data_in = testData5[4994];
@(posedge clk);
#1;data_in = testData5[4995];
@(posedge clk);
#1;data_in = testData5[4996];
@(posedge clk);
#1;data_in = testData5[4997];
@(posedge clk);
#1;data_in = testData5[4998];
@(posedge clk);
#1;data_in = testData5[4999];
@(posedge clk);
#1;data_in = testData5[5000];
@(posedge clk);
#1;data_in = testData5[5001];
@(posedge clk);
#1;data_in = testData5[5002];
@(posedge clk);
#1;data_in = testData5[5003];
@(posedge clk);
#1;data_in = testData5[5004];
@(posedge clk);
#1;data_in = testData5[5005];
@(posedge clk);
#1;data_in = testData5[5006];
@(posedge clk);
#1;data_in = testData5[5007];
@(posedge clk);
#1;data_in = testData5[5008];
@(posedge clk);
#1;data_in = testData5[5009];
@(posedge clk);
#1;data_in = testData5[5010];
@(posedge clk);
#1;data_in = testData5[5011];
@(posedge clk);
#1;data_in = testData5[5012];
@(posedge clk);
#1;data_in = testData5[5013];
@(posedge clk);
#1;data_in = testData5[5014];
@(posedge clk);
#1;data_in = testData5[5015];
@(posedge clk);
#1;data_in = testData5[5016];
@(posedge clk);
#1;data_in = testData5[5017];
@(posedge clk);
#1;data_in = testData5[5018];
@(posedge clk);
#1;data_in = testData5[5019];
@(posedge clk);
#1;data_in = testData5[5020];
@(posedge clk);
#1;data_in = testData5[5021];
@(posedge clk);
#1;data_in = testData5[5022];
@(posedge clk);
#1;data_in = testData5[5023];
@(posedge clk);
#1;data_in = testData5[5024];
@(posedge clk);
#1;data_in = testData5[5025];
@(posedge clk);
#1;data_in = testData5[5026];
@(posedge clk);
#1;data_in = testData5[5027];
@(posedge clk);
#1;data_in = testData5[5028];
@(posedge clk);
#1;data_in = testData5[5029];
@(posedge clk);
#1;data_in = testData5[5030];
@(posedge clk);
#1;data_in = testData5[5031];
@(posedge clk);
#1;data_in = testData5[5032];
@(posedge clk);
#1;data_in = testData5[5033];
@(posedge clk);
#1;data_in = testData5[5034];
@(posedge clk);
#1;data_in = testData5[5035];
@(posedge clk);
#1;data_in = testData5[5036];
@(posedge clk);
#1;data_in = testData5[5037];
@(posedge clk);
#1;data_in = testData5[5038];
@(posedge clk);
#1;data_in = testData5[5039];
@(posedge clk);
#1;data_in = testData5[5040];
@(posedge clk);
#1;data_in = testData5[5041];
@(posedge clk);
#1;data_in = testData5[5042];
@(posedge clk);
#1;data_in = testData5[5043];
@(posedge clk);
#1;data_in = testData5[5044];
@(posedge clk);
#1;data_in = testData5[5045];
@(posedge clk);
#1;data_in = testData5[5046];
@(posedge clk);
#1;data_in = testData5[5047];
@(posedge clk);
#1;data_in = testData5[5048];
@(posedge clk);
#1;data_in = testData5[5049];
@(posedge clk);
#1;data_in = testData5[5050];
@(posedge clk);
#1;data_in = testData5[5051];
@(posedge clk);
#1;data_in = testData5[5052];
@(posedge clk);
#1;data_in = testData5[5053];
@(posedge clk);
#1;data_in = testData5[5054];
@(posedge clk);
#1;data_in = testData5[5055];
@(posedge clk);
#1;data_in = testData5[5056];
@(posedge clk);
#1;data_in = testData5[5057];
@(posedge clk);
#1;data_in = testData5[5058];
@(posedge clk);
#1;data_in = testData5[5059];
@(posedge clk);
#1;data_in = testData5[5060];
@(posedge clk);
#1;data_in = testData5[5061];
@(posedge clk);
#1;data_in = testData5[5062];
@(posedge clk);
#1;data_in = testData5[5063];
@(posedge clk);
#1;data_in = testData5[5064];
@(posedge clk);
#1;data_in = testData5[5065];
@(posedge clk);
#1;data_in = testData5[5066];
@(posedge clk);
#1;data_in = testData5[5067];
@(posedge clk);
#1;data_in = testData5[5068];
@(posedge clk);
#1;data_in = testData5[5069];
@(posedge clk);
#1;data_in = testData5[5070];
@(posedge clk);
#1;data_in = testData5[5071];
@(posedge clk);
#1;data_in = testData5[5072];
@(posedge clk);
#1;data_in = testData5[5073];
@(posedge clk);
#1;data_in = testData5[5074];
@(posedge clk);
#1;data_in = testData5[5075];
@(posedge clk);
#1;data_in = testData5[5076];
@(posedge clk);
#1;data_in = testData5[5077];
@(posedge clk);
#1;data_in = testData5[5078];
@(posedge clk);
#1;data_in = testData5[5079];
@(posedge clk);
#1;data_in = testData5[5080];
@(posedge clk);
#1;data_in = testData5[5081];
@(posedge clk);
#1;data_in = testData5[5082];
@(posedge clk);
#1;data_in = testData5[5083];
@(posedge clk);
#1;data_in = testData5[5084];
@(posedge clk);
#1;data_in = testData5[5085];
@(posedge clk);
#1;data_in = testData5[5086];
@(posedge clk);
#1;data_in = testData5[5087];
@(posedge clk);
#1;data_in = testData5[5088];
@(posedge clk);
#1;data_in = testData5[5089];
@(posedge clk);
#1;data_in = testData5[5090];
@(posedge clk);
#1;data_in = testData5[5091];
@(posedge clk);
#1;data_in = testData5[5092];
@(posedge clk);
#1;data_in = testData5[5093];
@(posedge clk);
#1;data_in = testData5[5094];
@(posedge clk);
#1;data_in = testData5[5095];
@(posedge clk);
#1;data_in = testData5[5096];
@(posedge clk);
#1;data_in = testData5[5097];
@(posedge clk);
#1;data_in = testData5[5098];
@(posedge clk);
#1;data_in = testData5[5099];
@(posedge clk);
#1;data_in = testData5[5100];
@(posedge clk);
#1;data_in = testData5[5101];
@(posedge clk);
#1;data_in = testData5[5102];
@(posedge clk);
#1;data_in = testData5[5103];
@(posedge clk);
#1;data_in = testData5[5104];
@(posedge clk);
#1;data_in = testData5[5105];
@(posedge clk);
#1;data_in = testData5[5106];
@(posedge clk);
#1;data_in = testData5[5107];
@(posedge clk);
#1;data_in = testData5[5108];
@(posedge clk);
#1;data_in = testData5[5109];
@(posedge clk);
#1;data_in = testData5[5110];
@(posedge clk);
#1;data_in = testData5[5111];
@(posedge clk);
#1;data_in = testData5[5112];
@(posedge clk);
#1;data_in = testData5[5113];
@(posedge clk);
#1;data_in = testData5[5114];
@(posedge clk);
#1;data_in = testData5[5115];
@(posedge clk);
#1;data_in = testData5[5116];
@(posedge clk);
#1;data_in = testData5[5117];
@(posedge clk);
#1;data_in = testData5[5118];
@(posedge clk);
#1;data_in = testData5[5119];
@(posedge clk);
#1;data_in = testData5[5120];
@(posedge clk);
#1;data_in = testData5[5121];
@(posedge clk);
#1;data_in = testData5[5122];
@(posedge clk);
#1;data_in = testData5[5123];
@(posedge clk);
#1;data_in = testData5[5124];
@(posedge clk);
#1;data_in = testData5[5125];
@(posedge clk);
#1;data_in = testData5[5126];
@(posedge clk);
#1;data_in = testData5[5127];
@(posedge clk);
#1;data_in = testData5[5128];
@(posedge clk);
#1;data_in = testData5[5129];
@(posedge clk);
#1;data_in = testData5[5130];
@(posedge clk);
#1;data_in = testData5[5131];
@(posedge clk);
#1;data_in = testData5[5132];
@(posedge clk);
#1;data_in = testData5[5133];
@(posedge clk);
#1;data_in = testData5[5134];
@(posedge clk);
#1;data_in = testData5[5135];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[5136]; 
@(posedge clk);
#1;data_in = testData5[5137];
@(posedge clk);
#1;data_in = testData5[5138];
@(posedge clk);
#1;data_in = testData5[5139];
@(posedge clk);
#1;data_in = testData5[5140];
@(posedge clk);
#1;data_in = testData5[5141];
@(posedge clk);
#1;data_in = testData5[5142];
@(posedge clk);
#1;data_in = testData5[5143];
@(posedge clk);
#1;data_in = testData5[5144];
@(posedge clk);
#1;data_in = testData5[5145];
@(posedge clk);
#1;data_in = testData5[5146];
@(posedge clk);
#1;data_in = testData5[5147];
@(posedge clk);
#1;data_in = testData5[5148];
@(posedge clk);
#1;data_in = testData5[5149];
@(posedge clk);
#1;data_in = testData5[5150];
@(posedge clk);
#1;data_in = testData5[5151];
@(posedge clk);
#1;data_in = testData5[5152];
@(posedge clk);
#1;data_in = testData5[5153];
@(posedge clk);
#1;data_in = testData5[5154];
@(posedge clk);
#1;data_in = testData5[5155];
@(posedge clk);
#1;data_in = testData5[5156];
@(posedge clk);
#1;data_in = testData5[5157];
@(posedge clk);
#1;data_in = testData5[5158];
@(posedge clk);
#1;data_in = testData5[5159];
@(posedge clk);
#1;data_in = testData5[5160];
@(posedge clk);
#1;data_in = testData5[5161];
@(posedge clk);
#1;data_in = testData5[5162];
@(posedge clk);
#1;data_in = testData5[5163];
@(posedge clk);
#1;data_in = testData5[5164];
@(posedge clk);
#1;data_in = testData5[5165];
@(posedge clk);
#1;data_in = testData5[5166];
@(posedge clk);
#1;data_in = testData5[5167];
@(posedge clk);
#1;data_in = testData5[5168];
@(posedge clk);
#1;data_in = testData5[5169];
@(posedge clk);
#1;data_in = testData5[5170];
@(posedge clk);
#1;data_in = testData5[5171];
@(posedge clk);
#1;data_in = testData5[5172];
@(posedge clk);
#1;data_in = testData5[5173];
@(posedge clk);
#1;data_in = testData5[5174];
@(posedge clk);
#1;data_in = testData5[5175];
@(posedge clk);
#1;data_in = testData5[5176];
@(posedge clk);
#1;data_in = testData5[5177];
@(posedge clk);
#1;data_in = testData5[5178];
@(posedge clk);
#1;data_in = testData5[5179];
@(posedge clk);
#1;data_in = testData5[5180];
@(posedge clk);
#1;data_in = testData5[5181];
@(posedge clk);
#1;data_in = testData5[5182];
@(posedge clk);
#1;data_in = testData5[5183];
@(posedge clk);
#1;data_in = testData5[5184];
@(posedge clk);
#1;data_in = testData5[5185];
@(posedge clk);
#1;data_in = testData5[5186];
@(posedge clk);
#1;data_in = testData5[5187];
@(posedge clk);
#1;data_in = testData5[5188];
@(posedge clk);
#1;data_in = testData5[5189];
@(posedge clk);
#1;data_in = testData5[5190];
@(posedge clk);
#1;data_in = testData5[5191];
@(posedge clk);
#1;data_in = testData5[5192];
@(posedge clk);
#1;data_in = testData5[5193];
@(posedge clk);
#1;data_in = testData5[5194];
@(posedge clk);
#1;data_in = testData5[5195];
@(posedge clk);
#1;data_in = testData5[5196];
@(posedge clk);
#1;data_in = testData5[5197];
@(posedge clk);
#1;data_in = testData5[5198];
@(posedge clk);
#1;data_in = testData5[5199];
@(posedge clk);
#1;data_in = testData5[5200];
@(posedge clk);
#1;data_in = testData5[5201];
@(posedge clk);
#1;data_in = testData5[5202];
@(posedge clk);
#1;data_in = testData5[5203];
@(posedge clk);
#1;data_in = testData5[5204];
@(posedge clk);
#1;data_in = testData5[5205];
@(posedge clk);
#1;data_in = testData5[5206];
@(posedge clk);
#1;data_in = testData5[5207];
@(posedge clk);
#1;data_in = testData5[5208];
@(posedge clk);
#1;data_in = testData5[5209];
@(posedge clk);
#1;data_in = testData5[5210];
@(posedge clk);
#1;data_in = testData5[5211];
@(posedge clk);
#1;data_in = testData5[5212];
@(posedge clk);
#1;data_in = testData5[5213];
@(posedge clk);
#1;data_in = testData5[5214];
@(posedge clk);
#1;data_in = testData5[5215];
@(posedge clk);
#1;data_in = testData5[5216];
@(posedge clk);
#1;data_in = testData5[5217];
@(posedge clk);
#1;data_in = testData5[5218];
@(posedge clk);
#1;data_in = testData5[5219];
@(posedge clk);
#1;data_in = testData5[5220];
@(posedge clk);
#1;data_in = testData5[5221];
@(posedge clk);
#1;data_in = testData5[5222];
@(posedge clk);
#1;data_in = testData5[5223];
@(posedge clk);
#1;data_in = testData5[5224];
@(posedge clk);
#1;data_in = testData5[5225];
@(posedge clk);
#1;data_in = testData5[5226];
@(posedge clk);
#1;data_in = testData5[5227];
@(posedge clk);
#1;data_in = testData5[5228];
@(posedge clk);
#1;data_in = testData5[5229];
@(posedge clk);
#1;data_in = testData5[5230];
@(posedge clk);
#1;data_in = testData5[5231];
@(posedge clk);
#1;data_in = testData5[5232];
@(posedge clk);
#1;data_in = testData5[5233];
@(posedge clk);
#1;data_in = testData5[5234];
@(posedge clk);
#1;data_in = testData5[5235];
@(posedge clk);
#1;data_in = testData5[5236];
@(posedge clk);
#1;data_in = testData5[5237];
@(posedge clk);
#1;data_in = testData5[5238];
@(posedge clk);
#1;data_in = testData5[5239];
@(posedge clk);
#1;data_in = testData5[5240];
@(posedge clk);
#1;data_in = testData5[5241];
@(posedge clk);
#1;data_in = testData5[5242];
@(posedge clk);
#1;data_in = testData5[5243];
@(posedge clk);
#1;data_in = testData5[5244];
@(posedge clk);
#1;data_in = testData5[5245];
@(posedge clk);
#1;data_in = testData5[5246];
@(posedge clk);
#1;data_in = testData5[5247];
@(posedge clk);
#1;data_in = testData5[5248];
@(posedge clk);
#1;data_in = testData5[5249];
@(posedge clk);
#1;data_in = testData5[5250];
@(posedge clk);
#1;data_in = testData5[5251];
@(posedge clk);
#1;data_in = testData5[5252];
@(posedge clk);
#1;data_in = testData5[5253];
@(posedge clk);
#1;data_in = testData5[5254];
@(posedge clk);
#1;data_in = testData5[5255];
@(posedge clk);
#1;data_in = testData5[5256];
@(posedge clk);
#1;data_in = testData5[5257];
@(posedge clk);
#1;data_in = testData5[5258];
@(posedge clk);
#1;data_in = testData5[5259];
@(posedge clk);
#1;data_in = testData5[5260];
@(posedge clk);
#1;data_in = testData5[5261];
@(posedge clk);
#1;data_in = testData5[5262];
@(posedge clk);
#1;data_in = testData5[5263];
@(posedge clk);
#1;data_in = testData5[5264];
@(posedge clk);
#1;data_in = testData5[5265];
@(posedge clk);
#1;data_in = testData5[5266];
@(posedge clk);
#1;data_in = testData5[5267];
@(posedge clk);
#1;data_in = testData5[5268];
@(posedge clk);
#1;data_in = testData5[5269];
@(posedge clk);
#1;data_in = testData5[5270];
@(posedge clk);
#1;data_in = testData5[5271];
@(posedge clk);
#1;data_in = testData5[5272];
@(posedge clk);
#1;data_in = testData5[5273];
@(posedge clk);
#1;data_in = testData5[5274];
@(posedge clk);
#1;data_in = testData5[5275];
@(posedge clk);
#1;data_in = testData5[5276];
@(posedge clk);
#1;data_in = testData5[5277];
@(posedge clk);
#1;data_in = testData5[5278];
@(posedge clk);
#1;data_in = testData5[5279];
@(posedge clk);
#1;data_in = testData5[5280];
@(posedge clk);
#1;data_in = testData5[5281];
@(posedge clk);
#1;data_in = testData5[5282];
@(posedge clk);
#1;data_in = testData5[5283];
@(posedge clk);
#1;data_in = testData5[5284];
@(posedge clk);
#1;data_in = testData5[5285];
@(posedge clk);
#1;data_in = testData5[5286];
@(posedge clk);
#1;data_in = testData5[5287];
@(posedge clk);
#1;data_in = testData5[5288];
@(posedge clk);
#1;data_in = testData5[5289];
@(posedge clk);
#1;data_in = testData5[5290];
@(posedge clk);
#1;data_in = testData5[5291];
@(posedge clk);
#1;data_in = testData5[5292];
@(posedge clk);
#1;data_in = testData5[5293];
@(posedge clk);
#1;data_in = testData5[5294];
@(posedge clk);
#1;data_in = testData5[5295];
@(posedge clk);
#1;data_in = testData5[5296];
@(posedge clk);
#1;data_in = testData5[5297];
@(posedge clk);
#1;data_in = testData5[5298];
@(posedge clk);
#1;data_in = testData5[5299];
@(posedge clk);
#1;data_in = testData5[5300];
@(posedge clk);
#1;data_in = testData5[5301];
@(posedge clk);
#1;data_in = testData5[5302];
@(posedge clk);
#1;data_in = testData5[5303];
@(posedge clk);
#1;data_in = testData5[5304];
@(posedge clk);
#1;data_in = testData5[5305];
@(posedge clk);
#1;data_in = testData5[5306];
@(posedge clk);
#1;data_in = testData5[5307];
@(posedge clk);
#1;data_in = testData5[5308];
@(posedge clk);
#1;data_in = testData5[5309];
@(posedge clk);
#1;data_in = testData5[5310];
@(posedge clk);
#1;data_in = testData5[5311];
@(posedge clk);
#1;data_in = testData5[5312];
@(posedge clk);
#1;data_in = testData5[5313];
@(posedge clk);
#1;data_in = testData5[5314];
@(posedge clk);
#1;data_in = testData5[5315];
@(posedge clk);
#1;data_in = testData5[5316];
@(posedge clk);
#1;data_in = testData5[5317];
@(posedge clk);
#1;data_in = testData5[5318];
@(posedge clk);
#1;data_in = testData5[5319];
@(posedge clk);
#1;data_in = testData5[5320];
@(posedge clk);
#1;data_in = testData5[5321];
@(posedge clk);
#1;data_in = testData5[5322];
@(posedge clk);
#1;data_in = testData5[5323];
@(posedge clk);
#1;data_in = testData5[5324];
@(posedge clk);
#1;data_in = testData5[5325];
@(posedge clk);
#1;data_in = testData5[5326];
@(posedge clk);
#1;data_in = testData5[5327];
@(posedge clk);
#1;data_in = testData5[5328];
@(posedge clk);
#1;data_in = testData5[5329];
@(posedge clk);
#1;data_in = testData5[5330];
@(posedge clk);
#1;data_in = testData5[5331];
@(posedge clk);
#1;data_in = testData5[5332];
@(posedge clk);
#1;data_in = testData5[5333];
@(posedge clk);
#1;data_in = testData5[5334];
@(posedge clk);
#1;data_in = testData5[5335];
@(posedge clk);
#1;data_in = testData5[5336];
@(posedge clk);
#1;data_in = testData5[5337];
@(posedge clk);
#1;data_in = testData5[5338];
@(posedge clk);
#1;data_in = testData5[5339];
@(posedge clk);
#1;data_in = testData5[5340];
@(posedge clk);
#1;data_in = testData5[5341];
@(posedge clk);
#1;data_in = testData5[5342];
@(posedge clk);
#1;data_in = testData5[5343];
@(posedge clk);
#1;data_in = testData5[5344];
@(posedge clk);
#1;data_in = testData5[5345];
@(posedge clk);
#1;data_in = testData5[5346];
@(posedge clk);
#1;data_in = testData5[5347];
@(posedge clk);
#1;data_in = testData5[5348];
@(posedge clk);
#1;data_in = testData5[5349];
@(posedge clk);
#1;data_in = testData5[5350];
@(posedge clk);
#1;data_in = testData5[5351];
@(posedge clk);
#1;data_in = testData5[5352];
@(posedge clk);
#1;data_in = testData5[5353];
@(posedge clk);
#1;data_in = testData5[5354];
@(posedge clk);
#1;data_in = testData5[5355];
@(posedge clk);
#1;data_in = testData5[5356];
@(posedge clk);
#1;data_in = testData5[5357];
@(posedge clk);
#1;data_in = testData5[5358];
@(posedge clk);
#1;data_in = testData5[5359];
@(posedge clk);
#1;data_in = testData5[5360];
@(posedge clk);
#1;data_in = testData5[5361];
@(posedge clk);
#1;data_in = testData5[5362];
@(posedge clk);
#1;data_in = testData5[5363];
@(posedge clk);
#1;data_in = testData5[5364];
@(posedge clk);
#1;data_in = testData5[5365];
@(posedge clk);
#1;data_in = testData5[5366];
@(posedge clk);
#1;data_in = testData5[5367];
@(posedge clk);
#1;data_in = testData5[5368];
@(posedge clk);
#1;data_in = testData5[5369];
@(posedge clk);
#1;data_in = testData5[5370];
@(posedge clk);
#1;data_in = testData5[5371];
@(posedge clk);
#1;data_in = testData5[5372];
@(posedge clk);
#1;data_in = testData5[5373];
@(posedge clk);
#1;data_in = testData5[5374];
@(posedge clk);
#1;data_in = testData5[5375];
@(posedge clk);
#1;data_in = testData5[5376];
@(posedge clk);
#1;data_in = testData5[5377];
@(posedge clk);
#1;data_in = testData5[5378];
@(posedge clk);
#1;data_in = testData5[5379];
@(posedge clk);
#1;data_in = testData5[5380];
@(posedge clk);
#1;data_in = testData5[5381];
@(posedge clk);
#1;data_in = testData5[5382];
@(posedge clk);
#1;data_in = testData5[5383];
@(posedge clk);
#1;data_in = testData5[5384];
@(posedge clk);
#1;data_in = testData5[5385];
@(posedge clk);
#1;data_in = testData5[5386];
@(posedge clk);
#1;data_in = testData5[5387];
@(posedge clk);
#1;data_in = testData5[5388];
@(posedge clk);
#1;data_in = testData5[5389];
@(posedge clk);
#1;data_in = testData5[5390];
@(posedge clk);
#1;data_in = testData5[5391];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[5392]; 
@(posedge clk);
#1;data_in = testData5[5393];
@(posedge clk);
#1;data_in = testData5[5394];
@(posedge clk);
#1;data_in = testData5[5395];
@(posedge clk);
#1;data_in = testData5[5396];
@(posedge clk);
#1;data_in = testData5[5397];
@(posedge clk);
#1;data_in = testData5[5398];
@(posedge clk);
#1;data_in = testData5[5399];
@(posedge clk);
#1;data_in = testData5[5400];
@(posedge clk);
#1;data_in = testData5[5401];
@(posedge clk);
#1;data_in = testData5[5402];
@(posedge clk);
#1;data_in = testData5[5403];
@(posedge clk);
#1;data_in = testData5[5404];
@(posedge clk);
#1;data_in = testData5[5405];
@(posedge clk);
#1;data_in = testData5[5406];
@(posedge clk);
#1;data_in = testData5[5407];
@(posedge clk);
#1;data_in = testData5[5408];
@(posedge clk);
#1;data_in = testData5[5409];
@(posedge clk);
#1;data_in = testData5[5410];
@(posedge clk);
#1;data_in = testData5[5411];
@(posedge clk);
#1;data_in = testData5[5412];
@(posedge clk);
#1;data_in = testData5[5413];
@(posedge clk);
#1;data_in = testData5[5414];
@(posedge clk);
#1;data_in = testData5[5415];
@(posedge clk);
#1;data_in = testData5[5416];
@(posedge clk);
#1;data_in = testData5[5417];
@(posedge clk);
#1;data_in = testData5[5418];
@(posedge clk);
#1;data_in = testData5[5419];
@(posedge clk);
#1;data_in = testData5[5420];
@(posedge clk);
#1;data_in = testData5[5421];
@(posedge clk);
#1;data_in = testData5[5422];
@(posedge clk);
#1;data_in = testData5[5423];
@(posedge clk);
#1;data_in = testData5[5424];
@(posedge clk);
#1;data_in = testData5[5425];
@(posedge clk);
#1;data_in = testData5[5426];
@(posedge clk);
#1;data_in = testData5[5427];
@(posedge clk);
#1;data_in = testData5[5428];
@(posedge clk);
#1;data_in = testData5[5429];
@(posedge clk);
#1;data_in = testData5[5430];
@(posedge clk);
#1;data_in = testData5[5431];
@(posedge clk);
#1;data_in = testData5[5432];
@(posedge clk);
#1;data_in = testData5[5433];
@(posedge clk);
#1;data_in = testData5[5434];
@(posedge clk);
#1;data_in = testData5[5435];
@(posedge clk);
#1;data_in = testData5[5436];
@(posedge clk);
#1;data_in = testData5[5437];
@(posedge clk);
#1;data_in = testData5[5438];
@(posedge clk);
#1;data_in = testData5[5439];
@(posedge clk);
#1;data_in = testData5[5440];
@(posedge clk);
#1;data_in = testData5[5441];
@(posedge clk);
#1;data_in = testData5[5442];
@(posedge clk);
#1;data_in = testData5[5443];
@(posedge clk);
#1;data_in = testData5[5444];
@(posedge clk);
#1;data_in = testData5[5445];
@(posedge clk);
#1;data_in = testData5[5446];
@(posedge clk);
#1;data_in = testData5[5447];
@(posedge clk);
#1;data_in = testData5[5448];
@(posedge clk);
#1;data_in = testData5[5449];
@(posedge clk);
#1;data_in = testData5[5450];
@(posedge clk);
#1;data_in = testData5[5451];
@(posedge clk);
#1;data_in = testData5[5452];
@(posedge clk);
#1;data_in = testData5[5453];
@(posedge clk);
#1;data_in = testData5[5454];
@(posedge clk);
#1;data_in = testData5[5455];
@(posedge clk);
#1;data_in = testData5[5456];
@(posedge clk);
#1;data_in = testData5[5457];
@(posedge clk);
#1;data_in = testData5[5458];
@(posedge clk);
#1;data_in = testData5[5459];
@(posedge clk);
#1;data_in = testData5[5460];
@(posedge clk);
#1;data_in = testData5[5461];
@(posedge clk);
#1;data_in = testData5[5462];
@(posedge clk);
#1;data_in = testData5[5463];
@(posedge clk);
#1;data_in = testData5[5464];
@(posedge clk);
#1;data_in = testData5[5465];
@(posedge clk);
#1;data_in = testData5[5466];
@(posedge clk);
#1;data_in = testData5[5467];
@(posedge clk);
#1;data_in = testData5[5468];
@(posedge clk);
#1;data_in = testData5[5469];
@(posedge clk);
#1;data_in = testData5[5470];
@(posedge clk);
#1;data_in = testData5[5471];
@(posedge clk);
#1;data_in = testData5[5472];
@(posedge clk);
#1;data_in = testData5[5473];
@(posedge clk);
#1;data_in = testData5[5474];
@(posedge clk);
#1;data_in = testData5[5475];
@(posedge clk);
#1;data_in = testData5[5476];
@(posedge clk);
#1;data_in = testData5[5477];
@(posedge clk);
#1;data_in = testData5[5478];
@(posedge clk);
#1;data_in = testData5[5479];
@(posedge clk);
#1;data_in = testData5[5480];
@(posedge clk);
#1;data_in = testData5[5481];
@(posedge clk);
#1;data_in = testData5[5482];
@(posedge clk);
#1;data_in = testData5[5483];
@(posedge clk);
#1;data_in = testData5[5484];
@(posedge clk);
#1;data_in = testData5[5485];
@(posedge clk);
#1;data_in = testData5[5486];
@(posedge clk);
#1;data_in = testData5[5487];
@(posedge clk);
#1;data_in = testData5[5488];
@(posedge clk);
#1;data_in = testData5[5489];
@(posedge clk);
#1;data_in = testData5[5490];
@(posedge clk);
#1;data_in = testData5[5491];
@(posedge clk);
#1;data_in = testData5[5492];
@(posedge clk);
#1;data_in = testData5[5493];
@(posedge clk);
#1;data_in = testData5[5494];
@(posedge clk);
#1;data_in = testData5[5495];
@(posedge clk);
#1;data_in = testData5[5496];
@(posedge clk);
#1;data_in = testData5[5497];
@(posedge clk);
#1;data_in = testData5[5498];
@(posedge clk);
#1;data_in = testData5[5499];
@(posedge clk);
#1;data_in = testData5[5500];
@(posedge clk);
#1;data_in = testData5[5501];
@(posedge clk);
#1;data_in = testData5[5502];
@(posedge clk);
#1;data_in = testData5[5503];
@(posedge clk);
#1;data_in = testData5[5504];
@(posedge clk);
#1;data_in = testData5[5505];
@(posedge clk);
#1;data_in = testData5[5506];
@(posedge clk);
#1;data_in = testData5[5507];
@(posedge clk);
#1;data_in = testData5[5508];
@(posedge clk);
#1;data_in = testData5[5509];
@(posedge clk);
#1;data_in = testData5[5510];
@(posedge clk);
#1;data_in = testData5[5511];
@(posedge clk);
#1;data_in = testData5[5512];
@(posedge clk);
#1;data_in = testData5[5513];
@(posedge clk);
#1;data_in = testData5[5514];
@(posedge clk);
#1;data_in = testData5[5515];
@(posedge clk);
#1;data_in = testData5[5516];
@(posedge clk);
#1;data_in = testData5[5517];
@(posedge clk);
#1;data_in = testData5[5518];
@(posedge clk);
#1;data_in = testData5[5519];
@(posedge clk);
#1;data_in = testData5[5520];
@(posedge clk);
#1;data_in = testData5[5521];
@(posedge clk);
#1;data_in = testData5[5522];
@(posedge clk);
#1;data_in = testData5[5523];
@(posedge clk);
#1;data_in = testData5[5524];
@(posedge clk);
#1;data_in = testData5[5525];
@(posedge clk);
#1;data_in = testData5[5526];
@(posedge clk);
#1;data_in = testData5[5527];
@(posedge clk);
#1;data_in = testData5[5528];
@(posedge clk);
#1;data_in = testData5[5529];
@(posedge clk);
#1;data_in = testData5[5530];
@(posedge clk);
#1;data_in = testData5[5531];
@(posedge clk);
#1;data_in = testData5[5532];
@(posedge clk);
#1;data_in = testData5[5533];
@(posedge clk);
#1;data_in = testData5[5534];
@(posedge clk);
#1;data_in = testData5[5535];
@(posedge clk);
#1;data_in = testData5[5536];
@(posedge clk);
#1;data_in = testData5[5537];
@(posedge clk);
#1;data_in = testData5[5538];
@(posedge clk);
#1;data_in = testData5[5539];
@(posedge clk);
#1;data_in = testData5[5540];
@(posedge clk);
#1;data_in = testData5[5541];
@(posedge clk);
#1;data_in = testData5[5542];
@(posedge clk);
#1;data_in = testData5[5543];
@(posedge clk);
#1;data_in = testData5[5544];
@(posedge clk);
#1;data_in = testData5[5545];
@(posedge clk);
#1;data_in = testData5[5546];
@(posedge clk);
#1;data_in = testData5[5547];
@(posedge clk);
#1;data_in = testData5[5548];
@(posedge clk);
#1;data_in = testData5[5549];
@(posedge clk);
#1;data_in = testData5[5550];
@(posedge clk);
#1;data_in = testData5[5551];
@(posedge clk);
#1;data_in = testData5[5552];
@(posedge clk);
#1;data_in = testData5[5553];
@(posedge clk);
#1;data_in = testData5[5554];
@(posedge clk);
#1;data_in = testData5[5555];
@(posedge clk);
#1;data_in = testData5[5556];
@(posedge clk);
#1;data_in = testData5[5557];
@(posedge clk);
#1;data_in = testData5[5558];
@(posedge clk);
#1;data_in = testData5[5559];
@(posedge clk);
#1;data_in = testData5[5560];
@(posedge clk);
#1;data_in = testData5[5561];
@(posedge clk);
#1;data_in = testData5[5562];
@(posedge clk);
#1;data_in = testData5[5563];
@(posedge clk);
#1;data_in = testData5[5564];
@(posedge clk);
#1;data_in = testData5[5565];
@(posedge clk);
#1;data_in = testData5[5566];
@(posedge clk);
#1;data_in = testData5[5567];
@(posedge clk);
#1;data_in = testData5[5568];
@(posedge clk);
#1;data_in = testData5[5569];
@(posedge clk);
#1;data_in = testData5[5570];
@(posedge clk);
#1;data_in = testData5[5571];
@(posedge clk);
#1;data_in = testData5[5572];
@(posedge clk);
#1;data_in = testData5[5573];
@(posedge clk);
#1;data_in = testData5[5574];
@(posedge clk);
#1;data_in = testData5[5575];
@(posedge clk);
#1;data_in = testData5[5576];
@(posedge clk);
#1;data_in = testData5[5577];
@(posedge clk);
#1;data_in = testData5[5578];
@(posedge clk);
#1;data_in = testData5[5579];
@(posedge clk);
#1;data_in = testData5[5580];
@(posedge clk);
#1;data_in = testData5[5581];
@(posedge clk);
#1;data_in = testData5[5582];
@(posedge clk);
#1;data_in = testData5[5583];
@(posedge clk);
#1;data_in = testData5[5584];
@(posedge clk);
#1;data_in = testData5[5585];
@(posedge clk);
#1;data_in = testData5[5586];
@(posedge clk);
#1;data_in = testData5[5587];
@(posedge clk);
#1;data_in = testData5[5588];
@(posedge clk);
#1;data_in = testData5[5589];
@(posedge clk);
#1;data_in = testData5[5590];
@(posedge clk);
#1;data_in = testData5[5591];
@(posedge clk);
#1;data_in = testData5[5592];
@(posedge clk);
#1;data_in = testData5[5593];
@(posedge clk);
#1;data_in = testData5[5594];
@(posedge clk);
#1;data_in = testData5[5595];
@(posedge clk);
#1;data_in = testData5[5596];
@(posedge clk);
#1;data_in = testData5[5597];
@(posedge clk);
#1;data_in = testData5[5598];
@(posedge clk);
#1;data_in = testData5[5599];
@(posedge clk);
#1;data_in = testData5[5600];
@(posedge clk);
#1;data_in = testData5[5601];
@(posedge clk);
#1;data_in = testData5[5602];
@(posedge clk);
#1;data_in = testData5[5603];
@(posedge clk);
#1;data_in = testData5[5604];
@(posedge clk);
#1;data_in = testData5[5605];
@(posedge clk);
#1;data_in = testData5[5606];
@(posedge clk);
#1;data_in = testData5[5607];
@(posedge clk);
#1;data_in = testData5[5608];
@(posedge clk);
#1;data_in = testData5[5609];
@(posedge clk);
#1;data_in = testData5[5610];
@(posedge clk);
#1;data_in = testData5[5611];
@(posedge clk);
#1;data_in = testData5[5612];
@(posedge clk);
#1;data_in = testData5[5613];
@(posedge clk);
#1;data_in = testData5[5614];
@(posedge clk);
#1;data_in = testData5[5615];
@(posedge clk);
#1;data_in = testData5[5616];
@(posedge clk);
#1;data_in = testData5[5617];
@(posedge clk);
#1;data_in = testData5[5618];
@(posedge clk);
#1;data_in = testData5[5619];
@(posedge clk);
#1;data_in = testData5[5620];
@(posedge clk);
#1;data_in = testData5[5621];
@(posedge clk);
#1;data_in = testData5[5622];
@(posedge clk);
#1;data_in = testData5[5623];
@(posedge clk);
#1;data_in = testData5[5624];
@(posedge clk);
#1;data_in = testData5[5625];
@(posedge clk);
#1;data_in = testData5[5626];
@(posedge clk);
#1;data_in = testData5[5627];
@(posedge clk);
#1;data_in = testData5[5628];
@(posedge clk);
#1;data_in = testData5[5629];
@(posedge clk);
#1;data_in = testData5[5630];
@(posedge clk);
#1;data_in = testData5[5631];
@(posedge clk);
#1;data_in = testData5[5632];
@(posedge clk);
#1;data_in = testData5[5633];
@(posedge clk);
#1;data_in = testData5[5634];
@(posedge clk);
#1;data_in = testData5[5635];
@(posedge clk);
#1;data_in = testData5[5636];
@(posedge clk);
#1;data_in = testData5[5637];
@(posedge clk);
#1;data_in = testData5[5638];
@(posedge clk);
#1;data_in = testData5[5639];
@(posedge clk);
#1;data_in = testData5[5640];
@(posedge clk);
#1;data_in = testData5[5641];
@(posedge clk);
#1;data_in = testData5[5642];
@(posedge clk);
#1;data_in = testData5[5643];
@(posedge clk);
#1;data_in = testData5[5644];
@(posedge clk);
#1;data_in = testData5[5645];
@(posedge clk);
#1;data_in = testData5[5646];
@(posedge clk);
#1;data_in = testData5[5647];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[5648]; 
@(posedge clk);
#1;data_in = testData5[5649];
@(posedge clk);
#1;data_in = testData5[5650];
@(posedge clk);
#1;data_in = testData5[5651];
@(posedge clk);
#1;data_in = testData5[5652];
@(posedge clk);
#1;data_in = testData5[5653];
@(posedge clk);
#1;data_in = testData5[5654];
@(posedge clk);
#1;data_in = testData5[5655];
@(posedge clk);
#1;data_in = testData5[5656];
@(posedge clk);
#1;data_in = testData5[5657];
@(posedge clk);
#1;data_in = testData5[5658];
@(posedge clk);
#1;data_in = testData5[5659];
@(posedge clk);
#1;data_in = testData5[5660];
@(posedge clk);
#1;data_in = testData5[5661];
@(posedge clk);
#1;data_in = testData5[5662];
@(posedge clk);
#1;data_in = testData5[5663];
@(posedge clk);
#1;data_in = testData5[5664];
@(posedge clk);
#1;data_in = testData5[5665];
@(posedge clk);
#1;data_in = testData5[5666];
@(posedge clk);
#1;data_in = testData5[5667];
@(posedge clk);
#1;data_in = testData5[5668];
@(posedge clk);
#1;data_in = testData5[5669];
@(posedge clk);
#1;data_in = testData5[5670];
@(posedge clk);
#1;data_in = testData5[5671];
@(posedge clk);
#1;data_in = testData5[5672];
@(posedge clk);
#1;data_in = testData5[5673];
@(posedge clk);
#1;data_in = testData5[5674];
@(posedge clk);
#1;data_in = testData5[5675];
@(posedge clk);
#1;data_in = testData5[5676];
@(posedge clk);
#1;data_in = testData5[5677];
@(posedge clk);
#1;data_in = testData5[5678];
@(posedge clk);
#1;data_in = testData5[5679];
@(posedge clk);
#1;data_in = testData5[5680];
@(posedge clk);
#1;data_in = testData5[5681];
@(posedge clk);
#1;data_in = testData5[5682];
@(posedge clk);
#1;data_in = testData5[5683];
@(posedge clk);
#1;data_in = testData5[5684];
@(posedge clk);
#1;data_in = testData5[5685];
@(posedge clk);
#1;data_in = testData5[5686];
@(posedge clk);
#1;data_in = testData5[5687];
@(posedge clk);
#1;data_in = testData5[5688];
@(posedge clk);
#1;data_in = testData5[5689];
@(posedge clk);
#1;data_in = testData5[5690];
@(posedge clk);
#1;data_in = testData5[5691];
@(posedge clk);
#1;data_in = testData5[5692];
@(posedge clk);
#1;data_in = testData5[5693];
@(posedge clk);
#1;data_in = testData5[5694];
@(posedge clk);
#1;data_in = testData5[5695];
@(posedge clk);
#1;data_in = testData5[5696];
@(posedge clk);
#1;data_in = testData5[5697];
@(posedge clk);
#1;data_in = testData5[5698];
@(posedge clk);
#1;data_in = testData5[5699];
@(posedge clk);
#1;data_in = testData5[5700];
@(posedge clk);
#1;data_in = testData5[5701];
@(posedge clk);
#1;data_in = testData5[5702];
@(posedge clk);
#1;data_in = testData5[5703];
@(posedge clk);
#1;data_in = testData5[5704];
@(posedge clk);
#1;data_in = testData5[5705];
@(posedge clk);
#1;data_in = testData5[5706];
@(posedge clk);
#1;data_in = testData5[5707];
@(posedge clk);
#1;data_in = testData5[5708];
@(posedge clk);
#1;data_in = testData5[5709];
@(posedge clk);
#1;data_in = testData5[5710];
@(posedge clk);
#1;data_in = testData5[5711];
@(posedge clk);
#1;data_in = testData5[5712];
@(posedge clk);
#1;data_in = testData5[5713];
@(posedge clk);
#1;data_in = testData5[5714];
@(posedge clk);
#1;data_in = testData5[5715];
@(posedge clk);
#1;data_in = testData5[5716];
@(posedge clk);
#1;data_in = testData5[5717];
@(posedge clk);
#1;data_in = testData5[5718];
@(posedge clk);
#1;data_in = testData5[5719];
@(posedge clk);
#1;data_in = testData5[5720];
@(posedge clk);
#1;data_in = testData5[5721];
@(posedge clk);
#1;data_in = testData5[5722];
@(posedge clk);
#1;data_in = testData5[5723];
@(posedge clk);
#1;data_in = testData5[5724];
@(posedge clk);
#1;data_in = testData5[5725];
@(posedge clk);
#1;data_in = testData5[5726];
@(posedge clk);
#1;data_in = testData5[5727];
@(posedge clk);
#1;data_in = testData5[5728];
@(posedge clk);
#1;data_in = testData5[5729];
@(posedge clk);
#1;data_in = testData5[5730];
@(posedge clk);
#1;data_in = testData5[5731];
@(posedge clk);
#1;data_in = testData5[5732];
@(posedge clk);
#1;data_in = testData5[5733];
@(posedge clk);
#1;data_in = testData5[5734];
@(posedge clk);
#1;data_in = testData5[5735];
@(posedge clk);
#1;data_in = testData5[5736];
@(posedge clk);
#1;data_in = testData5[5737];
@(posedge clk);
#1;data_in = testData5[5738];
@(posedge clk);
#1;data_in = testData5[5739];
@(posedge clk);
#1;data_in = testData5[5740];
@(posedge clk);
#1;data_in = testData5[5741];
@(posedge clk);
#1;data_in = testData5[5742];
@(posedge clk);
#1;data_in = testData5[5743];
@(posedge clk);
#1;data_in = testData5[5744];
@(posedge clk);
#1;data_in = testData5[5745];
@(posedge clk);
#1;data_in = testData5[5746];
@(posedge clk);
#1;data_in = testData5[5747];
@(posedge clk);
#1;data_in = testData5[5748];
@(posedge clk);
#1;data_in = testData5[5749];
@(posedge clk);
#1;data_in = testData5[5750];
@(posedge clk);
#1;data_in = testData5[5751];
@(posedge clk);
#1;data_in = testData5[5752];
@(posedge clk);
#1;data_in = testData5[5753];
@(posedge clk);
#1;data_in = testData5[5754];
@(posedge clk);
#1;data_in = testData5[5755];
@(posedge clk);
#1;data_in = testData5[5756];
@(posedge clk);
#1;data_in = testData5[5757];
@(posedge clk);
#1;data_in = testData5[5758];
@(posedge clk);
#1;data_in = testData5[5759];
@(posedge clk);
#1;data_in = testData5[5760];
@(posedge clk);
#1;data_in = testData5[5761];
@(posedge clk);
#1;data_in = testData5[5762];
@(posedge clk);
#1;data_in = testData5[5763];
@(posedge clk);
#1;data_in = testData5[5764];
@(posedge clk);
#1;data_in = testData5[5765];
@(posedge clk);
#1;data_in = testData5[5766];
@(posedge clk);
#1;data_in = testData5[5767];
@(posedge clk);
#1;data_in = testData5[5768];
@(posedge clk);
#1;data_in = testData5[5769];
@(posedge clk);
#1;data_in = testData5[5770];
@(posedge clk);
#1;data_in = testData5[5771];
@(posedge clk);
#1;data_in = testData5[5772];
@(posedge clk);
#1;data_in = testData5[5773];
@(posedge clk);
#1;data_in = testData5[5774];
@(posedge clk);
#1;data_in = testData5[5775];
@(posedge clk);
#1;data_in = testData5[5776];
@(posedge clk);
#1;data_in = testData5[5777];
@(posedge clk);
#1;data_in = testData5[5778];
@(posedge clk);
#1;data_in = testData5[5779];
@(posedge clk);
#1;data_in = testData5[5780];
@(posedge clk);
#1;data_in = testData5[5781];
@(posedge clk);
#1;data_in = testData5[5782];
@(posedge clk);
#1;data_in = testData5[5783];
@(posedge clk);
#1;data_in = testData5[5784];
@(posedge clk);
#1;data_in = testData5[5785];
@(posedge clk);
#1;data_in = testData5[5786];
@(posedge clk);
#1;data_in = testData5[5787];
@(posedge clk);
#1;data_in = testData5[5788];
@(posedge clk);
#1;data_in = testData5[5789];
@(posedge clk);
#1;data_in = testData5[5790];
@(posedge clk);
#1;data_in = testData5[5791];
@(posedge clk);
#1;data_in = testData5[5792];
@(posedge clk);
#1;data_in = testData5[5793];
@(posedge clk);
#1;data_in = testData5[5794];
@(posedge clk);
#1;data_in = testData5[5795];
@(posedge clk);
#1;data_in = testData5[5796];
@(posedge clk);
#1;data_in = testData5[5797];
@(posedge clk);
#1;data_in = testData5[5798];
@(posedge clk);
#1;data_in = testData5[5799];
@(posedge clk);
#1;data_in = testData5[5800];
@(posedge clk);
#1;data_in = testData5[5801];
@(posedge clk);
#1;data_in = testData5[5802];
@(posedge clk);
#1;data_in = testData5[5803];
@(posedge clk);
#1;data_in = testData5[5804];
@(posedge clk);
#1;data_in = testData5[5805];
@(posedge clk);
#1;data_in = testData5[5806];
@(posedge clk);
#1;data_in = testData5[5807];
@(posedge clk);
#1;data_in = testData5[5808];
@(posedge clk);
#1;data_in = testData5[5809];
@(posedge clk);
#1;data_in = testData5[5810];
@(posedge clk);
#1;data_in = testData5[5811];
@(posedge clk);
#1;data_in = testData5[5812];
@(posedge clk);
#1;data_in = testData5[5813];
@(posedge clk);
#1;data_in = testData5[5814];
@(posedge clk);
#1;data_in = testData5[5815];
@(posedge clk);
#1;data_in = testData5[5816];
@(posedge clk);
#1;data_in = testData5[5817];
@(posedge clk);
#1;data_in = testData5[5818];
@(posedge clk);
#1;data_in = testData5[5819];
@(posedge clk);
#1;data_in = testData5[5820];
@(posedge clk);
#1;data_in = testData5[5821];
@(posedge clk);
#1;data_in = testData5[5822];
@(posedge clk);
#1;data_in = testData5[5823];
@(posedge clk);
#1;data_in = testData5[5824];
@(posedge clk);
#1;data_in = testData5[5825];
@(posedge clk);
#1;data_in = testData5[5826];
@(posedge clk);
#1;data_in = testData5[5827];
@(posedge clk);
#1;data_in = testData5[5828];
@(posedge clk);
#1;data_in = testData5[5829];
@(posedge clk);
#1;data_in = testData5[5830];
@(posedge clk);
#1;data_in = testData5[5831];
@(posedge clk);
#1;data_in = testData5[5832];
@(posedge clk);
#1;data_in = testData5[5833];
@(posedge clk);
#1;data_in = testData5[5834];
@(posedge clk);
#1;data_in = testData5[5835];
@(posedge clk);
#1;data_in = testData5[5836];
@(posedge clk);
#1;data_in = testData5[5837];
@(posedge clk);
#1;data_in = testData5[5838];
@(posedge clk);
#1;data_in = testData5[5839];
@(posedge clk);
#1;data_in = testData5[5840];
@(posedge clk);
#1;data_in = testData5[5841];
@(posedge clk);
#1;data_in = testData5[5842];
@(posedge clk);
#1;data_in = testData5[5843];
@(posedge clk);
#1;data_in = testData5[5844];
@(posedge clk);
#1;data_in = testData5[5845];
@(posedge clk);
#1;data_in = testData5[5846];
@(posedge clk);
#1;data_in = testData5[5847];
@(posedge clk);
#1;data_in = testData5[5848];
@(posedge clk);
#1;data_in = testData5[5849];
@(posedge clk);
#1;data_in = testData5[5850];
@(posedge clk);
#1;data_in = testData5[5851];
@(posedge clk);
#1;data_in = testData5[5852];
@(posedge clk);
#1;data_in = testData5[5853];
@(posedge clk);
#1;data_in = testData5[5854];
@(posedge clk);
#1;data_in = testData5[5855];
@(posedge clk);
#1;data_in = testData5[5856];
@(posedge clk);
#1;data_in = testData5[5857];
@(posedge clk);
#1;data_in = testData5[5858];
@(posedge clk);
#1;data_in = testData5[5859];
@(posedge clk);
#1;data_in = testData5[5860];
@(posedge clk);
#1;data_in = testData5[5861];
@(posedge clk);
#1;data_in = testData5[5862];
@(posedge clk);
#1;data_in = testData5[5863];
@(posedge clk);
#1;data_in = testData5[5864];
@(posedge clk);
#1;data_in = testData5[5865];
@(posedge clk);
#1;data_in = testData5[5866];
@(posedge clk);
#1;data_in = testData5[5867];
@(posedge clk);
#1;data_in = testData5[5868];
@(posedge clk);
#1;data_in = testData5[5869];
@(posedge clk);
#1;data_in = testData5[5870];
@(posedge clk);
#1;data_in = testData5[5871];
@(posedge clk);
#1;data_in = testData5[5872];
@(posedge clk);
#1;data_in = testData5[5873];
@(posedge clk);
#1;data_in = testData5[5874];
@(posedge clk);
#1;data_in = testData5[5875];
@(posedge clk);
#1;data_in = testData5[5876];
@(posedge clk);
#1;data_in = testData5[5877];
@(posedge clk);
#1;data_in = testData5[5878];
@(posedge clk);
#1;data_in = testData5[5879];
@(posedge clk);
#1;data_in = testData5[5880];
@(posedge clk);
#1;data_in = testData5[5881];
@(posedge clk);
#1;data_in = testData5[5882];
@(posedge clk);
#1;data_in = testData5[5883];
@(posedge clk);
#1;data_in = testData5[5884];
@(posedge clk);
#1;data_in = testData5[5885];
@(posedge clk);
#1;data_in = testData5[5886];
@(posedge clk);
#1;data_in = testData5[5887];
@(posedge clk);
#1;data_in = testData5[5888];
@(posedge clk);
#1;data_in = testData5[5889];
@(posedge clk);
#1;data_in = testData5[5890];
@(posedge clk);
#1;data_in = testData5[5891];
@(posedge clk);
#1;data_in = testData5[5892];
@(posedge clk);
#1;data_in = testData5[5893];
@(posedge clk);
#1;data_in = testData5[5894];
@(posedge clk);
#1;data_in = testData5[5895];
@(posedge clk);
#1;data_in = testData5[5896];
@(posedge clk);
#1;data_in = testData5[5897];
@(posedge clk);
#1;data_in = testData5[5898];
@(posedge clk);
#1;data_in = testData5[5899];
@(posedge clk);
#1;data_in = testData5[5900];
@(posedge clk);
#1;data_in = testData5[5901];
@(posedge clk);
#1;data_in = testData5[5902];
@(posedge clk);
#1;data_in = testData5[5903];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[5904]; 
@(posedge clk);
#1;data_in = testData5[5905];
@(posedge clk);
#1;data_in = testData5[5906];
@(posedge clk);
#1;data_in = testData5[5907];
@(posedge clk);
#1;data_in = testData5[5908];
@(posedge clk);
#1;data_in = testData5[5909];
@(posedge clk);
#1;data_in = testData5[5910];
@(posedge clk);
#1;data_in = testData5[5911];
@(posedge clk);
#1;data_in = testData5[5912];
@(posedge clk);
#1;data_in = testData5[5913];
@(posedge clk);
#1;data_in = testData5[5914];
@(posedge clk);
#1;data_in = testData5[5915];
@(posedge clk);
#1;data_in = testData5[5916];
@(posedge clk);
#1;data_in = testData5[5917];
@(posedge clk);
#1;data_in = testData5[5918];
@(posedge clk);
#1;data_in = testData5[5919];
@(posedge clk);
#1;data_in = testData5[5920];
@(posedge clk);
#1;data_in = testData5[5921];
@(posedge clk);
#1;data_in = testData5[5922];
@(posedge clk);
#1;data_in = testData5[5923];
@(posedge clk);
#1;data_in = testData5[5924];
@(posedge clk);
#1;data_in = testData5[5925];
@(posedge clk);
#1;data_in = testData5[5926];
@(posedge clk);
#1;data_in = testData5[5927];
@(posedge clk);
#1;data_in = testData5[5928];
@(posedge clk);
#1;data_in = testData5[5929];
@(posedge clk);
#1;data_in = testData5[5930];
@(posedge clk);
#1;data_in = testData5[5931];
@(posedge clk);
#1;data_in = testData5[5932];
@(posedge clk);
#1;data_in = testData5[5933];
@(posedge clk);
#1;data_in = testData5[5934];
@(posedge clk);
#1;data_in = testData5[5935];
@(posedge clk);
#1;data_in = testData5[5936];
@(posedge clk);
#1;data_in = testData5[5937];
@(posedge clk);
#1;data_in = testData5[5938];
@(posedge clk);
#1;data_in = testData5[5939];
@(posedge clk);
#1;data_in = testData5[5940];
@(posedge clk);
#1;data_in = testData5[5941];
@(posedge clk);
#1;data_in = testData5[5942];
@(posedge clk);
#1;data_in = testData5[5943];
@(posedge clk);
#1;data_in = testData5[5944];
@(posedge clk);
#1;data_in = testData5[5945];
@(posedge clk);
#1;data_in = testData5[5946];
@(posedge clk);
#1;data_in = testData5[5947];
@(posedge clk);
#1;data_in = testData5[5948];
@(posedge clk);
#1;data_in = testData5[5949];
@(posedge clk);
#1;data_in = testData5[5950];
@(posedge clk);
#1;data_in = testData5[5951];
@(posedge clk);
#1;data_in = testData5[5952];
@(posedge clk);
#1;data_in = testData5[5953];
@(posedge clk);
#1;data_in = testData5[5954];
@(posedge clk);
#1;data_in = testData5[5955];
@(posedge clk);
#1;data_in = testData5[5956];
@(posedge clk);
#1;data_in = testData5[5957];
@(posedge clk);
#1;data_in = testData5[5958];
@(posedge clk);
#1;data_in = testData5[5959];
@(posedge clk);
#1;data_in = testData5[5960];
@(posedge clk);
#1;data_in = testData5[5961];
@(posedge clk);
#1;data_in = testData5[5962];
@(posedge clk);
#1;data_in = testData5[5963];
@(posedge clk);
#1;data_in = testData5[5964];
@(posedge clk);
#1;data_in = testData5[5965];
@(posedge clk);
#1;data_in = testData5[5966];
@(posedge clk);
#1;data_in = testData5[5967];
@(posedge clk);
#1;data_in = testData5[5968];
@(posedge clk);
#1;data_in = testData5[5969];
@(posedge clk);
#1;data_in = testData5[5970];
@(posedge clk);
#1;data_in = testData5[5971];
@(posedge clk);
#1;data_in = testData5[5972];
@(posedge clk);
#1;data_in = testData5[5973];
@(posedge clk);
#1;data_in = testData5[5974];
@(posedge clk);
#1;data_in = testData5[5975];
@(posedge clk);
#1;data_in = testData5[5976];
@(posedge clk);
#1;data_in = testData5[5977];
@(posedge clk);
#1;data_in = testData5[5978];
@(posedge clk);
#1;data_in = testData5[5979];
@(posedge clk);
#1;data_in = testData5[5980];
@(posedge clk);
#1;data_in = testData5[5981];
@(posedge clk);
#1;data_in = testData5[5982];
@(posedge clk);
#1;data_in = testData5[5983];
@(posedge clk);
#1;data_in = testData5[5984];
@(posedge clk);
#1;data_in = testData5[5985];
@(posedge clk);
#1;data_in = testData5[5986];
@(posedge clk);
#1;data_in = testData5[5987];
@(posedge clk);
#1;data_in = testData5[5988];
@(posedge clk);
#1;data_in = testData5[5989];
@(posedge clk);
#1;data_in = testData5[5990];
@(posedge clk);
#1;data_in = testData5[5991];
@(posedge clk);
#1;data_in = testData5[5992];
@(posedge clk);
#1;data_in = testData5[5993];
@(posedge clk);
#1;data_in = testData5[5994];
@(posedge clk);
#1;data_in = testData5[5995];
@(posedge clk);
#1;data_in = testData5[5996];
@(posedge clk);
#1;data_in = testData5[5997];
@(posedge clk);
#1;data_in = testData5[5998];
@(posedge clk);
#1;data_in = testData5[5999];
@(posedge clk);
#1;data_in = testData5[6000];
@(posedge clk);
#1;data_in = testData5[6001];
@(posedge clk);
#1;data_in = testData5[6002];
@(posedge clk);
#1;data_in = testData5[6003];
@(posedge clk);
#1;data_in = testData5[6004];
@(posedge clk);
#1;data_in = testData5[6005];
@(posedge clk);
#1;data_in = testData5[6006];
@(posedge clk);
#1;data_in = testData5[6007];
@(posedge clk);
#1;data_in = testData5[6008];
@(posedge clk);
#1;data_in = testData5[6009];
@(posedge clk);
#1;data_in = testData5[6010];
@(posedge clk);
#1;data_in = testData5[6011];
@(posedge clk);
#1;data_in = testData5[6012];
@(posedge clk);
#1;data_in = testData5[6013];
@(posedge clk);
#1;data_in = testData5[6014];
@(posedge clk);
#1;data_in = testData5[6015];
@(posedge clk);
#1;data_in = testData5[6016];
@(posedge clk);
#1;data_in = testData5[6017];
@(posedge clk);
#1;data_in = testData5[6018];
@(posedge clk);
#1;data_in = testData5[6019];
@(posedge clk);
#1;data_in = testData5[6020];
@(posedge clk);
#1;data_in = testData5[6021];
@(posedge clk);
#1;data_in = testData5[6022];
@(posedge clk);
#1;data_in = testData5[6023];
@(posedge clk);
#1;data_in = testData5[6024];
@(posedge clk);
#1;data_in = testData5[6025];
@(posedge clk);
#1;data_in = testData5[6026];
@(posedge clk);
#1;data_in = testData5[6027];
@(posedge clk);
#1;data_in = testData5[6028];
@(posedge clk);
#1;data_in = testData5[6029];
@(posedge clk);
#1;data_in = testData5[6030];
@(posedge clk);
#1;data_in = testData5[6031];
@(posedge clk);
#1;data_in = testData5[6032];
@(posedge clk);
#1;data_in = testData5[6033];
@(posedge clk);
#1;data_in = testData5[6034];
@(posedge clk);
#1;data_in = testData5[6035];
@(posedge clk);
#1;data_in = testData5[6036];
@(posedge clk);
#1;data_in = testData5[6037];
@(posedge clk);
#1;data_in = testData5[6038];
@(posedge clk);
#1;data_in = testData5[6039];
@(posedge clk);
#1;data_in = testData5[6040];
@(posedge clk);
#1;data_in = testData5[6041];
@(posedge clk);
#1;data_in = testData5[6042];
@(posedge clk);
#1;data_in = testData5[6043];
@(posedge clk);
#1;data_in = testData5[6044];
@(posedge clk);
#1;data_in = testData5[6045];
@(posedge clk);
#1;data_in = testData5[6046];
@(posedge clk);
#1;data_in = testData5[6047];
@(posedge clk);
#1;data_in = testData5[6048];
@(posedge clk);
#1;data_in = testData5[6049];
@(posedge clk);
#1;data_in = testData5[6050];
@(posedge clk);
#1;data_in = testData5[6051];
@(posedge clk);
#1;data_in = testData5[6052];
@(posedge clk);
#1;data_in = testData5[6053];
@(posedge clk);
#1;data_in = testData5[6054];
@(posedge clk);
#1;data_in = testData5[6055];
@(posedge clk);
#1;data_in = testData5[6056];
@(posedge clk);
#1;data_in = testData5[6057];
@(posedge clk);
#1;data_in = testData5[6058];
@(posedge clk);
#1;data_in = testData5[6059];
@(posedge clk);
#1;data_in = testData5[6060];
@(posedge clk);
#1;data_in = testData5[6061];
@(posedge clk);
#1;data_in = testData5[6062];
@(posedge clk);
#1;data_in = testData5[6063];
@(posedge clk);
#1;data_in = testData5[6064];
@(posedge clk);
#1;data_in = testData5[6065];
@(posedge clk);
#1;data_in = testData5[6066];
@(posedge clk);
#1;data_in = testData5[6067];
@(posedge clk);
#1;data_in = testData5[6068];
@(posedge clk);
#1;data_in = testData5[6069];
@(posedge clk);
#1;data_in = testData5[6070];
@(posedge clk);
#1;data_in = testData5[6071];
@(posedge clk);
#1;data_in = testData5[6072];
@(posedge clk);
#1;data_in = testData5[6073];
@(posedge clk);
#1;data_in = testData5[6074];
@(posedge clk);
#1;data_in = testData5[6075];
@(posedge clk);
#1;data_in = testData5[6076];
@(posedge clk);
#1;data_in = testData5[6077];
@(posedge clk);
#1;data_in = testData5[6078];
@(posedge clk);
#1;data_in = testData5[6079];
@(posedge clk);
#1;data_in = testData5[6080];
@(posedge clk);
#1;data_in = testData5[6081];
@(posedge clk);
#1;data_in = testData5[6082];
@(posedge clk);
#1;data_in = testData5[6083];
@(posedge clk);
#1;data_in = testData5[6084];
@(posedge clk);
#1;data_in = testData5[6085];
@(posedge clk);
#1;data_in = testData5[6086];
@(posedge clk);
#1;data_in = testData5[6087];
@(posedge clk);
#1;data_in = testData5[6088];
@(posedge clk);
#1;data_in = testData5[6089];
@(posedge clk);
#1;data_in = testData5[6090];
@(posedge clk);
#1;data_in = testData5[6091];
@(posedge clk);
#1;data_in = testData5[6092];
@(posedge clk);
#1;data_in = testData5[6093];
@(posedge clk);
#1;data_in = testData5[6094];
@(posedge clk);
#1;data_in = testData5[6095];
@(posedge clk);
#1;data_in = testData5[6096];
@(posedge clk);
#1;data_in = testData5[6097];
@(posedge clk);
#1;data_in = testData5[6098];
@(posedge clk);
#1;data_in = testData5[6099];
@(posedge clk);
#1;data_in = testData5[6100];
@(posedge clk);
#1;data_in = testData5[6101];
@(posedge clk);
#1;data_in = testData5[6102];
@(posedge clk);
#1;data_in = testData5[6103];
@(posedge clk);
#1;data_in = testData5[6104];
@(posedge clk);
#1;data_in = testData5[6105];
@(posedge clk);
#1;data_in = testData5[6106];
@(posedge clk);
#1;data_in = testData5[6107];
@(posedge clk);
#1;data_in = testData5[6108];
@(posedge clk);
#1;data_in = testData5[6109];
@(posedge clk);
#1;data_in = testData5[6110];
@(posedge clk);
#1;data_in = testData5[6111];
@(posedge clk);
#1;data_in = testData5[6112];
@(posedge clk);
#1;data_in = testData5[6113];
@(posedge clk);
#1;data_in = testData5[6114];
@(posedge clk);
#1;data_in = testData5[6115];
@(posedge clk);
#1;data_in = testData5[6116];
@(posedge clk);
#1;data_in = testData5[6117];
@(posedge clk);
#1;data_in = testData5[6118];
@(posedge clk);
#1;data_in = testData5[6119];
@(posedge clk);
#1;data_in = testData5[6120];
@(posedge clk);
#1;data_in = testData5[6121];
@(posedge clk);
#1;data_in = testData5[6122];
@(posedge clk);
#1;data_in = testData5[6123];
@(posedge clk);
#1;data_in = testData5[6124];
@(posedge clk);
#1;data_in = testData5[6125];
@(posedge clk);
#1;data_in = testData5[6126];
@(posedge clk);
#1;data_in = testData5[6127];
@(posedge clk);
#1;data_in = testData5[6128];
@(posedge clk);
#1;data_in = testData5[6129];
@(posedge clk);
#1;data_in = testData5[6130];
@(posedge clk);
#1;data_in = testData5[6131];
@(posedge clk);
#1;data_in = testData5[6132];
@(posedge clk);
#1;data_in = testData5[6133];
@(posedge clk);
#1;data_in = testData5[6134];
@(posedge clk);
#1;data_in = testData5[6135];
@(posedge clk);
#1;data_in = testData5[6136];
@(posedge clk);
#1;data_in = testData5[6137];
@(posedge clk);
#1;data_in = testData5[6138];
@(posedge clk);
#1;data_in = testData5[6139];
@(posedge clk);
#1;data_in = testData5[6140];
@(posedge clk);
#1;data_in = testData5[6141];
@(posedge clk);
#1;data_in = testData5[6142];
@(posedge clk);
#1;data_in = testData5[6143];
@(posedge clk);
#1;data_in = testData5[6144];
@(posedge clk);
#1;data_in = testData5[6145];
@(posedge clk);
#1;data_in = testData5[6146];
@(posedge clk);
#1;data_in = testData5[6147];
@(posedge clk);
#1;data_in = testData5[6148];
@(posedge clk);
#1;data_in = testData5[6149];
@(posedge clk);
#1;data_in = testData5[6150];
@(posedge clk);
#1;data_in = testData5[6151];
@(posedge clk);
#1;data_in = testData5[6152];
@(posedge clk);
#1;data_in = testData5[6153];
@(posedge clk);
#1;data_in = testData5[6154];
@(posedge clk);
#1;data_in = testData5[6155];
@(posedge clk);
#1;data_in = testData5[6156];
@(posedge clk);
#1;data_in = testData5[6157];
@(posedge clk);
#1;data_in = testData5[6158];
@(posedge clk);
#1;data_in = testData5[6159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[6160]; 
@(posedge clk);
#1;data_in = testData5[6161];
@(posedge clk);
#1;data_in = testData5[6162];
@(posedge clk);
#1;data_in = testData5[6163];
@(posedge clk);
#1;data_in = testData5[6164];
@(posedge clk);
#1;data_in = testData5[6165];
@(posedge clk);
#1;data_in = testData5[6166];
@(posedge clk);
#1;data_in = testData5[6167];
@(posedge clk);
#1;data_in = testData5[6168];
@(posedge clk);
#1;data_in = testData5[6169];
@(posedge clk);
#1;data_in = testData5[6170];
@(posedge clk);
#1;data_in = testData5[6171];
@(posedge clk);
#1;data_in = testData5[6172];
@(posedge clk);
#1;data_in = testData5[6173];
@(posedge clk);
#1;data_in = testData5[6174];
@(posedge clk);
#1;data_in = testData5[6175];
@(posedge clk);
#1;data_in = testData5[6176];
@(posedge clk);
#1;data_in = testData5[6177];
@(posedge clk);
#1;data_in = testData5[6178];
@(posedge clk);
#1;data_in = testData5[6179];
@(posedge clk);
#1;data_in = testData5[6180];
@(posedge clk);
#1;data_in = testData5[6181];
@(posedge clk);
#1;data_in = testData5[6182];
@(posedge clk);
#1;data_in = testData5[6183];
@(posedge clk);
#1;data_in = testData5[6184];
@(posedge clk);
#1;data_in = testData5[6185];
@(posedge clk);
#1;data_in = testData5[6186];
@(posedge clk);
#1;data_in = testData5[6187];
@(posedge clk);
#1;data_in = testData5[6188];
@(posedge clk);
#1;data_in = testData5[6189];
@(posedge clk);
#1;data_in = testData5[6190];
@(posedge clk);
#1;data_in = testData5[6191];
@(posedge clk);
#1;data_in = testData5[6192];
@(posedge clk);
#1;data_in = testData5[6193];
@(posedge clk);
#1;data_in = testData5[6194];
@(posedge clk);
#1;data_in = testData5[6195];
@(posedge clk);
#1;data_in = testData5[6196];
@(posedge clk);
#1;data_in = testData5[6197];
@(posedge clk);
#1;data_in = testData5[6198];
@(posedge clk);
#1;data_in = testData5[6199];
@(posedge clk);
#1;data_in = testData5[6200];
@(posedge clk);
#1;data_in = testData5[6201];
@(posedge clk);
#1;data_in = testData5[6202];
@(posedge clk);
#1;data_in = testData5[6203];
@(posedge clk);
#1;data_in = testData5[6204];
@(posedge clk);
#1;data_in = testData5[6205];
@(posedge clk);
#1;data_in = testData5[6206];
@(posedge clk);
#1;data_in = testData5[6207];
@(posedge clk);
#1;data_in = testData5[6208];
@(posedge clk);
#1;data_in = testData5[6209];
@(posedge clk);
#1;data_in = testData5[6210];
@(posedge clk);
#1;data_in = testData5[6211];
@(posedge clk);
#1;data_in = testData5[6212];
@(posedge clk);
#1;data_in = testData5[6213];
@(posedge clk);
#1;data_in = testData5[6214];
@(posedge clk);
#1;data_in = testData5[6215];
@(posedge clk);
#1;data_in = testData5[6216];
@(posedge clk);
#1;data_in = testData5[6217];
@(posedge clk);
#1;data_in = testData5[6218];
@(posedge clk);
#1;data_in = testData5[6219];
@(posedge clk);
#1;data_in = testData5[6220];
@(posedge clk);
#1;data_in = testData5[6221];
@(posedge clk);
#1;data_in = testData5[6222];
@(posedge clk);
#1;data_in = testData5[6223];
@(posedge clk);
#1;data_in = testData5[6224];
@(posedge clk);
#1;data_in = testData5[6225];
@(posedge clk);
#1;data_in = testData5[6226];
@(posedge clk);
#1;data_in = testData5[6227];
@(posedge clk);
#1;data_in = testData5[6228];
@(posedge clk);
#1;data_in = testData5[6229];
@(posedge clk);
#1;data_in = testData5[6230];
@(posedge clk);
#1;data_in = testData5[6231];
@(posedge clk);
#1;data_in = testData5[6232];
@(posedge clk);
#1;data_in = testData5[6233];
@(posedge clk);
#1;data_in = testData5[6234];
@(posedge clk);
#1;data_in = testData5[6235];
@(posedge clk);
#1;data_in = testData5[6236];
@(posedge clk);
#1;data_in = testData5[6237];
@(posedge clk);
#1;data_in = testData5[6238];
@(posedge clk);
#1;data_in = testData5[6239];
@(posedge clk);
#1;data_in = testData5[6240];
@(posedge clk);
#1;data_in = testData5[6241];
@(posedge clk);
#1;data_in = testData5[6242];
@(posedge clk);
#1;data_in = testData5[6243];
@(posedge clk);
#1;data_in = testData5[6244];
@(posedge clk);
#1;data_in = testData5[6245];
@(posedge clk);
#1;data_in = testData5[6246];
@(posedge clk);
#1;data_in = testData5[6247];
@(posedge clk);
#1;data_in = testData5[6248];
@(posedge clk);
#1;data_in = testData5[6249];
@(posedge clk);
#1;data_in = testData5[6250];
@(posedge clk);
#1;data_in = testData5[6251];
@(posedge clk);
#1;data_in = testData5[6252];
@(posedge clk);
#1;data_in = testData5[6253];
@(posedge clk);
#1;data_in = testData5[6254];
@(posedge clk);
#1;data_in = testData5[6255];
@(posedge clk);
#1;data_in = testData5[6256];
@(posedge clk);
#1;data_in = testData5[6257];
@(posedge clk);
#1;data_in = testData5[6258];
@(posedge clk);
#1;data_in = testData5[6259];
@(posedge clk);
#1;data_in = testData5[6260];
@(posedge clk);
#1;data_in = testData5[6261];
@(posedge clk);
#1;data_in = testData5[6262];
@(posedge clk);
#1;data_in = testData5[6263];
@(posedge clk);
#1;data_in = testData5[6264];
@(posedge clk);
#1;data_in = testData5[6265];
@(posedge clk);
#1;data_in = testData5[6266];
@(posedge clk);
#1;data_in = testData5[6267];
@(posedge clk);
#1;data_in = testData5[6268];
@(posedge clk);
#1;data_in = testData5[6269];
@(posedge clk);
#1;data_in = testData5[6270];
@(posedge clk);
#1;data_in = testData5[6271];
@(posedge clk);
#1;data_in = testData5[6272];
@(posedge clk);
#1;data_in = testData5[6273];
@(posedge clk);
#1;data_in = testData5[6274];
@(posedge clk);
#1;data_in = testData5[6275];
@(posedge clk);
#1;data_in = testData5[6276];
@(posedge clk);
#1;data_in = testData5[6277];
@(posedge clk);
#1;data_in = testData5[6278];
@(posedge clk);
#1;data_in = testData5[6279];
@(posedge clk);
#1;data_in = testData5[6280];
@(posedge clk);
#1;data_in = testData5[6281];
@(posedge clk);
#1;data_in = testData5[6282];
@(posedge clk);
#1;data_in = testData5[6283];
@(posedge clk);
#1;data_in = testData5[6284];
@(posedge clk);
#1;data_in = testData5[6285];
@(posedge clk);
#1;data_in = testData5[6286];
@(posedge clk);
#1;data_in = testData5[6287];
@(posedge clk);
#1;data_in = testData5[6288];
@(posedge clk);
#1;data_in = testData5[6289];
@(posedge clk);
#1;data_in = testData5[6290];
@(posedge clk);
#1;data_in = testData5[6291];
@(posedge clk);
#1;data_in = testData5[6292];
@(posedge clk);
#1;data_in = testData5[6293];
@(posedge clk);
#1;data_in = testData5[6294];
@(posedge clk);
#1;data_in = testData5[6295];
@(posedge clk);
#1;data_in = testData5[6296];
@(posedge clk);
#1;data_in = testData5[6297];
@(posedge clk);
#1;data_in = testData5[6298];
@(posedge clk);
#1;data_in = testData5[6299];
@(posedge clk);
#1;data_in = testData5[6300];
@(posedge clk);
#1;data_in = testData5[6301];
@(posedge clk);
#1;data_in = testData5[6302];
@(posedge clk);
#1;data_in = testData5[6303];
@(posedge clk);
#1;data_in = testData5[6304];
@(posedge clk);
#1;data_in = testData5[6305];
@(posedge clk);
#1;data_in = testData5[6306];
@(posedge clk);
#1;data_in = testData5[6307];
@(posedge clk);
#1;data_in = testData5[6308];
@(posedge clk);
#1;data_in = testData5[6309];
@(posedge clk);
#1;data_in = testData5[6310];
@(posedge clk);
#1;data_in = testData5[6311];
@(posedge clk);
#1;data_in = testData5[6312];
@(posedge clk);
#1;data_in = testData5[6313];
@(posedge clk);
#1;data_in = testData5[6314];
@(posedge clk);
#1;data_in = testData5[6315];
@(posedge clk);
#1;data_in = testData5[6316];
@(posedge clk);
#1;data_in = testData5[6317];
@(posedge clk);
#1;data_in = testData5[6318];
@(posedge clk);
#1;data_in = testData5[6319];
@(posedge clk);
#1;data_in = testData5[6320];
@(posedge clk);
#1;data_in = testData5[6321];
@(posedge clk);
#1;data_in = testData5[6322];
@(posedge clk);
#1;data_in = testData5[6323];
@(posedge clk);
#1;data_in = testData5[6324];
@(posedge clk);
#1;data_in = testData5[6325];
@(posedge clk);
#1;data_in = testData5[6326];
@(posedge clk);
#1;data_in = testData5[6327];
@(posedge clk);
#1;data_in = testData5[6328];
@(posedge clk);
#1;data_in = testData5[6329];
@(posedge clk);
#1;data_in = testData5[6330];
@(posedge clk);
#1;data_in = testData5[6331];
@(posedge clk);
#1;data_in = testData5[6332];
@(posedge clk);
#1;data_in = testData5[6333];
@(posedge clk);
#1;data_in = testData5[6334];
@(posedge clk);
#1;data_in = testData5[6335];
@(posedge clk);
#1;data_in = testData5[6336];
@(posedge clk);
#1;data_in = testData5[6337];
@(posedge clk);
#1;data_in = testData5[6338];
@(posedge clk);
#1;data_in = testData5[6339];
@(posedge clk);
#1;data_in = testData5[6340];
@(posedge clk);
#1;data_in = testData5[6341];
@(posedge clk);
#1;data_in = testData5[6342];
@(posedge clk);
#1;data_in = testData5[6343];
@(posedge clk);
#1;data_in = testData5[6344];
@(posedge clk);
#1;data_in = testData5[6345];
@(posedge clk);
#1;data_in = testData5[6346];
@(posedge clk);
#1;data_in = testData5[6347];
@(posedge clk);
#1;data_in = testData5[6348];
@(posedge clk);
#1;data_in = testData5[6349];
@(posedge clk);
#1;data_in = testData5[6350];
@(posedge clk);
#1;data_in = testData5[6351];
@(posedge clk);
#1;data_in = testData5[6352];
@(posedge clk);
#1;data_in = testData5[6353];
@(posedge clk);
#1;data_in = testData5[6354];
@(posedge clk);
#1;data_in = testData5[6355];
@(posedge clk);
#1;data_in = testData5[6356];
@(posedge clk);
#1;data_in = testData5[6357];
@(posedge clk);
#1;data_in = testData5[6358];
@(posedge clk);
#1;data_in = testData5[6359];
@(posedge clk);
#1;data_in = testData5[6360];
@(posedge clk);
#1;data_in = testData5[6361];
@(posedge clk);
#1;data_in = testData5[6362];
@(posedge clk);
#1;data_in = testData5[6363];
@(posedge clk);
#1;data_in = testData5[6364];
@(posedge clk);
#1;data_in = testData5[6365];
@(posedge clk);
#1;data_in = testData5[6366];
@(posedge clk);
#1;data_in = testData5[6367];
@(posedge clk);
#1;data_in = testData5[6368];
@(posedge clk);
#1;data_in = testData5[6369];
@(posedge clk);
#1;data_in = testData5[6370];
@(posedge clk);
#1;data_in = testData5[6371];
@(posedge clk);
#1;data_in = testData5[6372];
@(posedge clk);
#1;data_in = testData5[6373];
@(posedge clk);
#1;data_in = testData5[6374];
@(posedge clk);
#1;data_in = testData5[6375];
@(posedge clk);
#1;data_in = testData5[6376];
@(posedge clk);
#1;data_in = testData5[6377];
@(posedge clk);
#1;data_in = testData5[6378];
@(posedge clk);
#1;data_in = testData5[6379];
@(posedge clk);
#1;data_in = testData5[6380];
@(posedge clk);
#1;data_in = testData5[6381];
@(posedge clk);
#1;data_in = testData5[6382];
@(posedge clk);
#1;data_in = testData5[6383];
@(posedge clk);
#1;data_in = testData5[6384];
@(posedge clk);
#1;data_in = testData5[6385];
@(posedge clk);
#1;data_in = testData5[6386];
@(posedge clk);
#1;data_in = testData5[6387];
@(posedge clk);
#1;data_in = testData5[6388];
@(posedge clk);
#1;data_in = testData5[6389];
@(posedge clk);
#1;data_in = testData5[6390];
@(posedge clk);
#1;data_in = testData5[6391];
@(posedge clk);
#1;data_in = testData5[6392];
@(posedge clk);
#1;data_in = testData5[6393];
@(posedge clk);
#1;data_in = testData5[6394];
@(posedge clk);
#1;data_in = testData5[6395];
@(posedge clk);
#1;data_in = testData5[6396];
@(posedge clk);
#1;data_in = testData5[6397];
@(posedge clk);
#1;data_in = testData5[6398];
@(posedge clk);
#1;data_in = testData5[6399];
@(posedge clk);
#1;data_in = testData5[6400];
@(posedge clk);
#1;data_in = testData5[6401];
@(posedge clk);
#1;data_in = testData5[6402];
@(posedge clk);
#1;data_in = testData5[6403];
@(posedge clk);
#1;data_in = testData5[6404];
@(posedge clk);
#1;data_in = testData5[6405];
@(posedge clk);
#1;data_in = testData5[6406];
@(posedge clk);
#1;data_in = testData5[6407];
@(posedge clk);
#1;data_in = testData5[6408];
@(posedge clk);
#1;data_in = testData5[6409];
@(posedge clk);
#1;data_in = testData5[6410];
@(posedge clk);
#1;data_in = testData5[6411];
@(posedge clk);
#1;data_in = testData5[6412];
@(posedge clk);
#1;data_in = testData5[6413];
@(posedge clk);
#1;data_in = testData5[6414];
@(posedge clk);
#1;data_in = testData5[6415];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[6416]; 
@(posedge clk);
#1;data_in = testData5[6417];
@(posedge clk);
#1;data_in = testData5[6418];
@(posedge clk);
#1;data_in = testData5[6419];
@(posedge clk);
#1;data_in = testData5[6420];
@(posedge clk);
#1;data_in = testData5[6421];
@(posedge clk);
#1;data_in = testData5[6422];
@(posedge clk);
#1;data_in = testData5[6423];
@(posedge clk);
#1;data_in = testData5[6424];
@(posedge clk);
#1;data_in = testData5[6425];
@(posedge clk);
#1;data_in = testData5[6426];
@(posedge clk);
#1;data_in = testData5[6427];
@(posedge clk);
#1;data_in = testData5[6428];
@(posedge clk);
#1;data_in = testData5[6429];
@(posedge clk);
#1;data_in = testData5[6430];
@(posedge clk);
#1;data_in = testData5[6431];
@(posedge clk);
#1;data_in = testData5[6432];
@(posedge clk);
#1;data_in = testData5[6433];
@(posedge clk);
#1;data_in = testData5[6434];
@(posedge clk);
#1;data_in = testData5[6435];
@(posedge clk);
#1;data_in = testData5[6436];
@(posedge clk);
#1;data_in = testData5[6437];
@(posedge clk);
#1;data_in = testData5[6438];
@(posedge clk);
#1;data_in = testData5[6439];
@(posedge clk);
#1;data_in = testData5[6440];
@(posedge clk);
#1;data_in = testData5[6441];
@(posedge clk);
#1;data_in = testData5[6442];
@(posedge clk);
#1;data_in = testData5[6443];
@(posedge clk);
#1;data_in = testData5[6444];
@(posedge clk);
#1;data_in = testData5[6445];
@(posedge clk);
#1;data_in = testData5[6446];
@(posedge clk);
#1;data_in = testData5[6447];
@(posedge clk);
#1;data_in = testData5[6448];
@(posedge clk);
#1;data_in = testData5[6449];
@(posedge clk);
#1;data_in = testData5[6450];
@(posedge clk);
#1;data_in = testData5[6451];
@(posedge clk);
#1;data_in = testData5[6452];
@(posedge clk);
#1;data_in = testData5[6453];
@(posedge clk);
#1;data_in = testData5[6454];
@(posedge clk);
#1;data_in = testData5[6455];
@(posedge clk);
#1;data_in = testData5[6456];
@(posedge clk);
#1;data_in = testData5[6457];
@(posedge clk);
#1;data_in = testData5[6458];
@(posedge clk);
#1;data_in = testData5[6459];
@(posedge clk);
#1;data_in = testData5[6460];
@(posedge clk);
#1;data_in = testData5[6461];
@(posedge clk);
#1;data_in = testData5[6462];
@(posedge clk);
#1;data_in = testData5[6463];
@(posedge clk);
#1;data_in = testData5[6464];
@(posedge clk);
#1;data_in = testData5[6465];
@(posedge clk);
#1;data_in = testData5[6466];
@(posedge clk);
#1;data_in = testData5[6467];
@(posedge clk);
#1;data_in = testData5[6468];
@(posedge clk);
#1;data_in = testData5[6469];
@(posedge clk);
#1;data_in = testData5[6470];
@(posedge clk);
#1;data_in = testData5[6471];
@(posedge clk);
#1;data_in = testData5[6472];
@(posedge clk);
#1;data_in = testData5[6473];
@(posedge clk);
#1;data_in = testData5[6474];
@(posedge clk);
#1;data_in = testData5[6475];
@(posedge clk);
#1;data_in = testData5[6476];
@(posedge clk);
#1;data_in = testData5[6477];
@(posedge clk);
#1;data_in = testData5[6478];
@(posedge clk);
#1;data_in = testData5[6479];
@(posedge clk);
#1;data_in = testData5[6480];
@(posedge clk);
#1;data_in = testData5[6481];
@(posedge clk);
#1;data_in = testData5[6482];
@(posedge clk);
#1;data_in = testData5[6483];
@(posedge clk);
#1;data_in = testData5[6484];
@(posedge clk);
#1;data_in = testData5[6485];
@(posedge clk);
#1;data_in = testData5[6486];
@(posedge clk);
#1;data_in = testData5[6487];
@(posedge clk);
#1;data_in = testData5[6488];
@(posedge clk);
#1;data_in = testData5[6489];
@(posedge clk);
#1;data_in = testData5[6490];
@(posedge clk);
#1;data_in = testData5[6491];
@(posedge clk);
#1;data_in = testData5[6492];
@(posedge clk);
#1;data_in = testData5[6493];
@(posedge clk);
#1;data_in = testData5[6494];
@(posedge clk);
#1;data_in = testData5[6495];
@(posedge clk);
#1;data_in = testData5[6496];
@(posedge clk);
#1;data_in = testData5[6497];
@(posedge clk);
#1;data_in = testData5[6498];
@(posedge clk);
#1;data_in = testData5[6499];
@(posedge clk);
#1;data_in = testData5[6500];
@(posedge clk);
#1;data_in = testData5[6501];
@(posedge clk);
#1;data_in = testData5[6502];
@(posedge clk);
#1;data_in = testData5[6503];
@(posedge clk);
#1;data_in = testData5[6504];
@(posedge clk);
#1;data_in = testData5[6505];
@(posedge clk);
#1;data_in = testData5[6506];
@(posedge clk);
#1;data_in = testData5[6507];
@(posedge clk);
#1;data_in = testData5[6508];
@(posedge clk);
#1;data_in = testData5[6509];
@(posedge clk);
#1;data_in = testData5[6510];
@(posedge clk);
#1;data_in = testData5[6511];
@(posedge clk);
#1;data_in = testData5[6512];
@(posedge clk);
#1;data_in = testData5[6513];
@(posedge clk);
#1;data_in = testData5[6514];
@(posedge clk);
#1;data_in = testData5[6515];
@(posedge clk);
#1;data_in = testData5[6516];
@(posedge clk);
#1;data_in = testData5[6517];
@(posedge clk);
#1;data_in = testData5[6518];
@(posedge clk);
#1;data_in = testData5[6519];
@(posedge clk);
#1;data_in = testData5[6520];
@(posedge clk);
#1;data_in = testData5[6521];
@(posedge clk);
#1;data_in = testData5[6522];
@(posedge clk);
#1;data_in = testData5[6523];
@(posedge clk);
#1;data_in = testData5[6524];
@(posedge clk);
#1;data_in = testData5[6525];
@(posedge clk);
#1;data_in = testData5[6526];
@(posedge clk);
#1;data_in = testData5[6527];
@(posedge clk);
#1;data_in = testData5[6528];
@(posedge clk);
#1;data_in = testData5[6529];
@(posedge clk);
#1;data_in = testData5[6530];
@(posedge clk);
#1;data_in = testData5[6531];
@(posedge clk);
#1;data_in = testData5[6532];
@(posedge clk);
#1;data_in = testData5[6533];
@(posedge clk);
#1;data_in = testData5[6534];
@(posedge clk);
#1;data_in = testData5[6535];
@(posedge clk);
#1;data_in = testData5[6536];
@(posedge clk);
#1;data_in = testData5[6537];
@(posedge clk);
#1;data_in = testData5[6538];
@(posedge clk);
#1;data_in = testData5[6539];
@(posedge clk);
#1;data_in = testData5[6540];
@(posedge clk);
#1;data_in = testData5[6541];
@(posedge clk);
#1;data_in = testData5[6542];
@(posedge clk);
#1;data_in = testData5[6543];
@(posedge clk);
#1;data_in = testData5[6544];
@(posedge clk);
#1;data_in = testData5[6545];
@(posedge clk);
#1;data_in = testData5[6546];
@(posedge clk);
#1;data_in = testData5[6547];
@(posedge clk);
#1;data_in = testData5[6548];
@(posedge clk);
#1;data_in = testData5[6549];
@(posedge clk);
#1;data_in = testData5[6550];
@(posedge clk);
#1;data_in = testData5[6551];
@(posedge clk);
#1;data_in = testData5[6552];
@(posedge clk);
#1;data_in = testData5[6553];
@(posedge clk);
#1;data_in = testData5[6554];
@(posedge clk);
#1;data_in = testData5[6555];
@(posedge clk);
#1;data_in = testData5[6556];
@(posedge clk);
#1;data_in = testData5[6557];
@(posedge clk);
#1;data_in = testData5[6558];
@(posedge clk);
#1;data_in = testData5[6559];
@(posedge clk);
#1;data_in = testData5[6560];
@(posedge clk);
#1;data_in = testData5[6561];
@(posedge clk);
#1;data_in = testData5[6562];
@(posedge clk);
#1;data_in = testData5[6563];
@(posedge clk);
#1;data_in = testData5[6564];
@(posedge clk);
#1;data_in = testData5[6565];
@(posedge clk);
#1;data_in = testData5[6566];
@(posedge clk);
#1;data_in = testData5[6567];
@(posedge clk);
#1;data_in = testData5[6568];
@(posedge clk);
#1;data_in = testData5[6569];
@(posedge clk);
#1;data_in = testData5[6570];
@(posedge clk);
#1;data_in = testData5[6571];
@(posedge clk);
#1;data_in = testData5[6572];
@(posedge clk);
#1;data_in = testData5[6573];
@(posedge clk);
#1;data_in = testData5[6574];
@(posedge clk);
#1;data_in = testData5[6575];
@(posedge clk);
#1;data_in = testData5[6576];
@(posedge clk);
#1;data_in = testData5[6577];
@(posedge clk);
#1;data_in = testData5[6578];
@(posedge clk);
#1;data_in = testData5[6579];
@(posedge clk);
#1;data_in = testData5[6580];
@(posedge clk);
#1;data_in = testData5[6581];
@(posedge clk);
#1;data_in = testData5[6582];
@(posedge clk);
#1;data_in = testData5[6583];
@(posedge clk);
#1;data_in = testData5[6584];
@(posedge clk);
#1;data_in = testData5[6585];
@(posedge clk);
#1;data_in = testData5[6586];
@(posedge clk);
#1;data_in = testData5[6587];
@(posedge clk);
#1;data_in = testData5[6588];
@(posedge clk);
#1;data_in = testData5[6589];
@(posedge clk);
#1;data_in = testData5[6590];
@(posedge clk);
#1;data_in = testData5[6591];
@(posedge clk);
#1;data_in = testData5[6592];
@(posedge clk);
#1;data_in = testData5[6593];
@(posedge clk);
#1;data_in = testData5[6594];
@(posedge clk);
#1;data_in = testData5[6595];
@(posedge clk);
#1;data_in = testData5[6596];
@(posedge clk);
#1;data_in = testData5[6597];
@(posedge clk);
#1;data_in = testData5[6598];
@(posedge clk);
#1;data_in = testData5[6599];
@(posedge clk);
#1;data_in = testData5[6600];
@(posedge clk);
#1;data_in = testData5[6601];
@(posedge clk);
#1;data_in = testData5[6602];
@(posedge clk);
#1;data_in = testData5[6603];
@(posedge clk);
#1;data_in = testData5[6604];
@(posedge clk);
#1;data_in = testData5[6605];
@(posedge clk);
#1;data_in = testData5[6606];
@(posedge clk);
#1;data_in = testData5[6607];
@(posedge clk);
#1;data_in = testData5[6608];
@(posedge clk);
#1;data_in = testData5[6609];
@(posedge clk);
#1;data_in = testData5[6610];
@(posedge clk);
#1;data_in = testData5[6611];
@(posedge clk);
#1;data_in = testData5[6612];
@(posedge clk);
#1;data_in = testData5[6613];
@(posedge clk);
#1;data_in = testData5[6614];
@(posedge clk);
#1;data_in = testData5[6615];
@(posedge clk);
#1;data_in = testData5[6616];
@(posedge clk);
#1;data_in = testData5[6617];
@(posedge clk);
#1;data_in = testData5[6618];
@(posedge clk);
#1;data_in = testData5[6619];
@(posedge clk);
#1;data_in = testData5[6620];
@(posedge clk);
#1;data_in = testData5[6621];
@(posedge clk);
#1;data_in = testData5[6622];
@(posedge clk);
#1;data_in = testData5[6623];
@(posedge clk);
#1;data_in = testData5[6624];
@(posedge clk);
#1;data_in = testData5[6625];
@(posedge clk);
#1;data_in = testData5[6626];
@(posedge clk);
#1;data_in = testData5[6627];
@(posedge clk);
#1;data_in = testData5[6628];
@(posedge clk);
#1;data_in = testData5[6629];
@(posedge clk);
#1;data_in = testData5[6630];
@(posedge clk);
#1;data_in = testData5[6631];
@(posedge clk);
#1;data_in = testData5[6632];
@(posedge clk);
#1;data_in = testData5[6633];
@(posedge clk);
#1;data_in = testData5[6634];
@(posedge clk);
#1;data_in = testData5[6635];
@(posedge clk);
#1;data_in = testData5[6636];
@(posedge clk);
#1;data_in = testData5[6637];
@(posedge clk);
#1;data_in = testData5[6638];
@(posedge clk);
#1;data_in = testData5[6639];
@(posedge clk);
#1;data_in = testData5[6640];
@(posedge clk);
#1;data_in = testData5[6641];
@(posedge clk);
#1;data_in = testData5[6642];
@(posedge clk);
#1;data_in = testData5[6643];
@(posedge clk);
#1;data_in = testData5[6644];
@(posedge clk);
#1;data_in = testData5[6645];
@(posedge clk);
#1;data_in = testData5[6646];
@(posedge clk);
#1;data_in = testData5[6647];
@(posedge clk);
#1;data_in = testData5[6648];
@(posedge clk);
#1;data_in = testData5[6649];
@(posedge clk);
#1;data_in = testData5[6650];
@(posedge clk);
#1;data_in = testData5[6651];
@(posedge clk);
#1;data_in = testData5[6652];
@(posedge clk);
#1;data_in = testData5[6653];
@(posedge clk);
#1;data_in = testData5[6654];
@(posedge clk);
#1;data_in = testData5[6655];
@(posedge clk);
#1;data_in = testData5[6656];
@(posedge clk);
#1;data_in = testData5[6657];
@(posedge clk);
#1;data_in = testData5[6658];
@(posedge clk);
#1;data_in = testData5[6659];
@(posedge clk);
#1;data_in = testData5[6660];
@(posedge clk);
#1;data_in = testData5[6661];
@(posedge clk);
#1;data_in = testData5[6662];
@(posedge clk);
#1;data_in = testData5[6663];
@(posedge clk);
#1;data_in = testData5[6664];
@(posedge clk);
#1;data_in = testData5[6665];
@(posedge clk);
#1;data_in = testData5[6666];
@(posedge clk);
#1;data_in = testData5[6667];
@(posedge clk);
#1;data_in = testData5[6668];
@(posedge clk);
#1;data_in = testData5[6669];
@(posedge clk);
#1;data_in = testData5[6670];
@(posedge clk);
#1;data_in = testData5[6671];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[6672]; 
@(posedge clk);
#1;data_in = testData5[6673];
@(posedge clk);
#1;data_in = testData5[6674];
@(posedge clk);
#1;data_in = testData5[6675];
@(posedge clk);
#1;data_in = testData5[6676];
@(posedge clk);
#1;data_in = testData5[6677];
@(posedge clk);
#1;data_in = testData5[6678];
@(posedge clk);
#1;data_in = testData5[6679];
@(posedge clk);
#1;data_in = testData5[6680];
@(posedge clk);
#1;data_in = testData5[6681];
@(posedge clk);
#1;data_in = testData5[6682];
@(posedge clk);
#1;data_in = testData5[6683];
@(posedge clk);
#1;data_in = testData5[6684];
@(posedge clk);
#1;data_in = testData5[6685];
@(posedge clk);
#1;data_in = testData5[6686];
@(posedge clk);
#1;data_in = testData5[6687];
@(posedge clk);
#1;data_in = testData5[6688];
@(posedge clk);
#1;data_in = testData5[6689];
@(posedge clk);
#1;data_in = testData5[6690];
@(posedge clk);
#1;data_in = testData5[6691];
@(posedge clk);
#1;data_in = testData5[6692];
@(posedge clk);
#1;data_in = testData5[6693];
@(posedge clk);
#1;data_in = testData5[6694];
@(posedge clk);
#1;data_in = testData5[6695];
@(posedge clk);
#1;data_in = testData5[6696];
@(posedge clk);
#1;data_in = testData5[6697];
@(posedge clk);
#1;data_in = testData5[6698];
@(posedge clk);
#1;data_in = testData5[6699];
@(posedge clk);
#1;data_in = testData5[6700];
@(posedge clk);
#1;data_in = testData5[6701];
@(posedge clk);
#1;data_in = testData5[6702];
@(posedge clk);
#1;data_in = testData5[6703];
@(posedge clk);
#1;data_in = testData5[6704];
@(posedge clk);
#1;data_in = testData5[6705];
@(posedge clk);
#1;data_in = testData5[6706];
@(posedge clk);
#1;data_in = testData5[6707];
@(posedge clk);
#1;data_in = testData5[6708];
@(posedge clk);
#1;data_in = testData5[6709];
@(posedge clk);
#1;data_in = testData5[6710];
@(posedge clk);
#1;data_in = testData5[6711];
@(posedge clk);
#1;data_in = testData5[6712];
@(posedge clk);
#1;data_in = testData5[6713];
@(posedge clk);
#1;data_in = testData5[6714];
@(posedge clk);
#1;data_in = testData5[6715];
@(posedge clk);
#1;data_in = testData5[6716];
@(posedge clk);
#1;data_in = testData5[6717];
@(posedge clk);
#1;data_in = testData5[6718];
@(posedge clk);
#1;data_in = testData5[6719];
@(posedge clk);
#1;data_in = testData5[6720];
@(posedge clk);
#1;data_in = testData5[6721];
@(posedge clk);
#1;data_in = testData5[6722];
@(posedge clk);
#1;data_in = testData5[6723];
@(posedge clk);
#1;data_in = testData5[6724];
@(posedge clk);
#1;data_in = testData5[6725];
@(posedge clk);
#1;data_in = testData5[6726];
@(posedge clk);
#1;data_in = testData5[6727];
@(posedge clk);
#1;data_in = testData5[6728];
@(posedge clk);
#1;data_in = testData5[6729];
@(posedge clk);
#1;data_in = testData5[6730];
@(posedge clk);
#1;data_in = testData5[6731];
@(posedge clk);
#1;data_in = testData5[6732];
@(posedge clk);
#1;data_in = testData5[6733];
@(posedge clk);
#1;data_in = testData5[6734];
@(posedge clk);
#1;data_in = testData5[6735];
@(posedge clk);
#1;data_in = testData5[6736];
@(posedge clk);
#1;data_in = testData5[6737];
@(posedge clk);
#1;data_in = testData5[6738];
@(posedge clk);
#1;data_in = testData5[6739];
@(posedge clk);
#1;data_in = testData5[6740];
@(posedge clk);
#1;data_in = testData5[6741];
@(posedge clk);
#1;data_in = testData5[6742];
@(posedge clk);
#1;data_in = testData5[6743];
@(posedge clk);
#1;data_in = testData5[6744];
@(posedge clk);
#1;data_in = testData5[6745];
@(posedge clk);
#1;data_in = testData5[6746];
@(posedge clk);
#1;data_in = testData5[6747];
@(posedge clk);
#1;data_in = testData5[6748];
@(posedge clk);
#1;data_in = testData5[6749];
@(posedge clk);
#1;data_in = testData5[6750];
@(posedge clk);
#1;data_in = testData5[6751];
@(posedge clk);
#1;data_in = testData5[6752];
@(posedge clk);
#1;data_in = testData5[6753];
@(posedge clk);
#1;data_in = testData5[6754];
@(posedge clk);
#1;data_in = testData5[6755];
@(posedge clk);
#1;data_in = testData5[6756];
@(posedge clk);
#1;data_in = testData5[6757];
@(posedge clk);
#1;data_in = testData5[6758];
@(posedge clk);
#1;data_in = testData5[6759];
@(posedge clk);
#1;data_in = testData5[6760];
@(posedge clk);
#1;data_in = testData5[6761];
@(posedge clk);
#1;data_in = testData5[6762];
@(posedge clk);
#1;data_in = testData5[6763];
@(posedge clk);
#1;data_in = testData5[6764];
@(posedge clk);
#1;data_in = testData5[6765];
@(posedge clk);
#1;data_in = testData5[6766];
@(posedge clk);
#1;data_in = testData5[6767];
@(posedge clk);
#1;data_in = testData5[6768];
@(posedge clk);
#1;data_in = testData5[6769];
@(posedge clk);
#1;data_in = testData5[6770];
@(posedge clk);
#1;data_in = testData5[6771];
@(posedge clk);
#1;data_in = testData5[6772];
@(posedge clk);
#1;data_in = testData5[6773];
@(posedge clk);
#1;data_in = testData5[6774];
@(posedge clk);
#1;data_in = testData5[6775];
@(posedge clk);
#1;data_in = testData5[6776];
@(posedge clk);
#1;data_in = testData5[6777];
@(posedge clk);
#1;data_in = testData5[6778];
@(posedge clk);
#1;data_in = testData5[6779];
@(posedge clk);
#1;data_in = testData5[6780];
@(posedge clk);
#1;data_in = testData5[6781];
@(posedge clk);
#1;data_in = testData5[6782];
@(posedge clk);
#1;data_in = testData5[6783];
@(posedge clk);
#1;data_in = testData5[6784];
@(posedge clk);
#1;data_in = testData5[6785];
@(posedge clk);
#1;data_in = testData5[6786];
@(posedge clk);
#1;data_in = testData5[6787];
@(posedge clk);
#1;data_in = testData5[6788];
@(posedge clk);
#1;data_in = testData5[6789];
@(posedge clk);
#1;data_in = testData5[6790];
@(posedge clk);
#1;data_in = testData5[6791];
@(posedge clk);
#1;data_in = testData5[6792];
@(posedge clk);
#1;data_in = testData5[6793];
@(posedge clk);
#1;data_in = testData5[6794];
@(posedge clk);
#1;data_in = testData5[6795];
@(posedge clk);
#1;data_in = testData5[6796];
@(posedge clk);
#1;data_in = testData5[6797];
@(posedge clk);
#1;data_in = testData5[6798];
@(posedge clk);
#1;data_in = testData5[6799];
@(posedge clk);
#1;data_in = testData5[6800];
@(posedge clk);
#1;data_in = testData5[6801];
@(posedge clk);
#1;data_in = testData5[6802];
@(posedge clk);
#1;data_in = testData5[6803];
@(posedge clk);
#1;data_in = testData5[6804];
@(posedge clk);
#1;data_in = testData5[6805];
@(posedge clk);
#1;data_in = testData5[6806];
@(posedge clk);
#1;data_in = testData5[6807];
@(posedge clk);
#1;data_in = testData5[6808];
@(posedge clk);
#1;data_in = testData5[6809];
@(posedge clk);
#1;data_in = testData5[6810];
@(posedge clk);
#1;data_in = testData5[6811];
@(posedge clk);
#1;data_in = testData5[6812];
@(posedge clk);
#1;data_in = testData5[6813];
@(posedge clk);
#1;data_in = testData5[6814];
@(posedge clk);
#1;data_in = testData5[6815];
@(posedge clk);
#1;data_in = testData5[6816];
@(posedge clk);
#1;data_in = testData5[6817];
@(posedge clk);
#1;data_in = testData5[6818];
@(posedge clk);
#1;data_in = testData5[6819];
@(posedge clk);
#1;data_in = testData5[6820];
@(posedge clk);
#1;data_in = testData5[6821];
@(posedge clk);
#1;data_in = testData5[6822];
@(posedge clk);
#1;data_in = testData5[6823];
@(posedge clk);
#1;data_in = testData5[6824];
@(posedge clk);
#1;data_in = testData5[6825];
@(posedge clk);
#1;data_in = testData5[6826];
@(posedge clk);
#1;data_in = testData5[6827];
@(posedge clk);
#1;data_in = testData5[6828];
@(posedge clk);
#1;data_in = testData5[6829];
@(posedge clk);
#1;data_in = testData5[6830];
@(posedge clk);
#1;data_in = testData5[6831];
@(posedge clk);
#1;data_in = testData5[6832];
@(posedge clk);
#1;data_in = testData5[6833];
@(posedge clk);
#1;data_in = testData5[6834];
@(posedge clk);
#1;data_in = testData5[6835];
@(posedge clk);
#1;data_in = testData5[6836];
@(posedge clk);
#1;data_in = testData5[6837];
@(posedge clk);
#1;data_in = testData5[6838];
@(posedge clk);
#1;data_in = testData5[6839];
@(posedge clk);
#1;data_in = testData5[6840];
@(posedge clk);
#1;data_in = testData5[6841];
@(posedge clk);
#1;data_in = testData5[6842];
@(posedge clk);
#1;data_in = testData5[6843];
@(posedge clk);
#1;data_in = testData5[6844];
@(posedge clk);
#1;data_in = testData5[6845];
@(posedge clk);
#1;data_in = testData5[6846];
@(posedge clk);
#1;data_in = testData5[6847];
@(posedge clk);
#1;data_in = testData5[6848];
@(posedge clk);
#1;data_in = testData5[6849];
@(posedge clk);
#1;data_in = testData5[6850];
@(posedge clk);
#1;data_in = testData5[6851];
@(posedge clk);
#1;data_in = testData5[6852];
@(posedge clk);
#1;data_in = testData5[6853];
@(posedge clk);
#1;data_in = testData5[6854];
@(posedge clk);
#1;data_in = testData5[6855];
@(posedge clk);
#1;data_in = testData5[6856];
@(posedge clk);
#1;data_in = testData5[6857];
@(posedge clk);
#1;data_in = testData5[6858];
@(posedge clk);
#1;data_in = testData5[6859];
@(posedge clk);
#1;data_in = testData5[6860];
@(posedge clk);
#1;data_in = testData5[6861];
@(posedge clk);
#1;data_in = testData5[6862];
@(posedge clk);
#1;data_in = testData5[6863];
@(posedge clk);
#1;data_in = testData5[6864];
@(posedge clk);
#1;data_in = testData5[6865];
@(posedge clk);
#1;data_in = testData5[6866];
@(posedge clk);
#1;data_in = testData5[6867];
@(posedge clk);
#1;data_in = testData5[6868];
@(posedge clk);
#1;data_in = testData5[6869];
@(posedge clk);
#1;data_in = testData5[6870];
@(posedge clk);
#1;data_in = testData5[6871];
@(posedge clk);
#1;data_in = testData5[6872];
@(posedge clk);
#1;data_in = testData5[6873];
@(posedge clk);
#1;data_in = testData5[6874];
@(posedge clk);
#1;data_in = testData5[6875];
@(posedge clk);
#1;data_in = testData5[6876];
@(posedge clk);
#1;data_in = testData5[6877];
@(posedge clk);
#1;data_in = testData5[6878];
@(posedge clk);
#1;data_in = testData5[6879];
@(posedge clk);
#1;data_in = testData5[6880];
@(posedge clk);
#1;data_in = testData5[6881];
@(posedge clk);
#1;data_in = testData5[6882];
@(posedge clk);
#1;data_in = testData5[6883];
@(posedge clk);
#1;data_in = testData5[6884];
@(posedge clk);
#1;data_in = testData5[6885];
@(posedge clk);
#1;data_in = testData5[6886];
@(posedge clk);
#1;data_in = testData5[6887];
@(posedge clk);
#1;data_in = testData5[6888];
@(posedge clk);
#1;data_in = testData5[6889];
@(posedge clk);
#1;data_in = testData5[6890];
@(posedge clk);
#1;data_in = testData5[6891];
@(posedge clk);
#1;data_in = testData5[6892];
@(posedge clk);
#1;data_in = testData5[6893];
@(posedge clk);
#1;data_in = testData5[6894];
@(posedge clk);
#1;data_in = testData5[6895];
@(posedge clk);
#1;data_in = testData5[6896];
@(posedge clk);
#1;data_in = testData5[6897];
@(posedge clk);
#1;data_in = testData5[6898];
@(posedge clk);
#1;data_in = testData5[6899];
@(posedge clk);
#1;data_in = testData5[6900];
@(posedge clk);
#1;data_in = testData5[6901];
@(posedge clk);
#1;data_in = testData5[6902];
@(posedge clk);
#1;data_in = testData5[6903];
@(posedge clk);
#1;data_in = testData5[6904];
@(posedge clk);
#1;data_in = testData5[6905];
@(posedge clk);
#1;data_in = testData5[6906];
@(posedge clk);
#1;data_in = testData5[6907];
@(posedge clk);
#1;data_in = testData5[6908];
@(posedge clk);
#1;data_in = testData5[6909];
@(posedge clk);
#1;data_in = testData5[6910];
@(posedge clk);
#1;data_in = testData5[6911];
@(posedge clk);
#1;data_in = testData5[6912];
@(posedge clk);
#1;data_in = testData5[6913];
@(posedge clk);
#1;data_in = testData5[6914];
@(posedge clk);
#1;data_in = testData5[6915];
@(posedge clk);
#1;data_in = testData5[6916];
@(posedge clk);
#1;data_in = testData5[6917];
@(posedge clk);
#1;data_in = testData5[6918];
@(posedge clk);
#1;data_in = testData5[6919];
@(posedge clk);
#1;data_in = testData5[6920];
@(posedge clk);
#1;data_in = testData5[6921];
@(posedge clk);
#1;data_in = testData5[6922];
@(posedge clk);
#1;data_in = testData5[6923];
@(posedge clk);
#1;data_in = testData5[6924];
@(posedge clk);
#1;data_in = testData5[6925];
@(posedge clk);
#1;data_in = testData5[6926];
@(posedge clk);
#1;data_in = testData5[6927];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[6928]; 
@(posedge clk);
#1;data_in = testData5[6929];
@(posedge clk);
#1;data_in = testData5[6930];
@(posedge clk);
#1;data_in = testData5[6931];
@(posedge clk);
#1;data_in = testData5[6932];
@(posedge clk);
#1;data_in = testData5[6933];
@(posedge clk);
#1;data_in = testData5[6934];
@(posedge clk);
#1;data_in = testData5[6935];
@(posedge clk);
#1;data_in = testData5[6936];
@(posedge clk);
#1;data_in = testData5[6937];
@(posedge clk);
#1;data_in = testData5[6938];
@(posedge clk);
#1;data_in = testData5[6939];
@(posedge clk);
#1;data_in = testData5[6940];
@(posedge clk);
#1;data_in = testData5[6941];
@(posedge clk);
#1;data_in = testData5[6942];
@(posedge clk);
#1;data_in = testData5[6943];
@(posedge clk);
#1;data_in = testData5[6944];
@(posedge clk);
#1;data_in = testData5[6945];
@(posedge clk);
#1;data_in = testData5[6946];
@(posedge clk);
#1;data_in = testData5[6947];
@(posedge clk);
#1;data_in = testData5[6948];
@(posedge clk);
#1;data_in = testData5[6949];
@(posedge clk);
#1;data_in = testData5[6950];
@(posedge clk);
#1;data_in = testData5[6951];
@(posedge clk);
#1;data_in = testData5[6952];
@(posedge clk);
#1;data_in = testData5[6953];
@(posedge clk);
#1;data_in = testData5[6954];
@(posedge clk);
#1;data_in = testData5[6955];
@(posedge clk);
#1;data_in = testData5[6956];
@(posedge clk);
#1;data_in = testData5[6957];
@(posedge clk);
#1;data_in = testData5[6958];
@(posedge clk);
#1;data_in = testData5[6959];
@(posedge clk);
#1;data_in = testData5[6960];
@(posedge clk);
#1;data_in = testData5[6961];
@(posedge clk);
#1;data_in = testData5[6962];
@(posedge clk);
#1;data_in = testData5[6963];
@(posedge clk);
#1;data_in = testData5[6964];
@(posedge clk);
#1;data_in = testData5[6965];
@(posedge clk);
#1;data_in = testData5[6966];
@(posedge clk);
#1;data_in = testData5[6967];
@(posedge clk);
#1;data_in = testData5[6968];
@(posedge clk);
#1;data_in = testData5[6969];
@(posedge clk);
#1;data_in = testData5[6970];
@(posedge clk);
#1;data_in = testData5[6971];
@(posedge clk);
#1;data_in = testData5[6972];
@(posedge clk);
#1;data_in = testData5[6973];
@(posedge clk);
#1;data_in = testData5[6974];
@(posedge clk);
#1;data_in = testData5[6975];
@(posedge clk);
#1;data_in = testData5[6976];
@(posedge clk);
#1;data_in = testData5[6977];
@(posedge clk);
#1;data_in = testData5[6978];
@(posedge clk);
#1;data_in = testData5[6979];
@(posedge clk);
#1;data_in = testData5[6980];
@(posedge clk);
#1;data_in = testData5[6981];
@(posedge clk);
#1;data_in = testData5[6982];
@(posedge clk);
#1;data_in = testData5[6983];
@(posedge clk);
#1;data_in = testData5[6984];
@(posedge clk);
#1;data_in = testData5[6985];
@(posedge clk);
#1;data_in = testData5[6986];
@(posedge clk);
#1;data_in = testData5[6987];
@(posedge clk);
#1;data_in = testData5[6988];
@(posedge clk);
#1;data_in = testData5[6989];
@(posedge clk);
#1;data_in = testData5[6990];
@(posedge clk);
#1;data_in = testData5[6991];
@(posedge clk);
#1;data_in = testData5[6992];
@(posedge clk);
#1;data_in = testData5[6993];
@(posedge clk);
#1;data_in = testData5[6994];
@(posedge clk);
#1;data_in = testData5[6995];
@(posedge clk);
#1;data_in = testData5[6996];
@(posedge clk);
#1;data_in = testData5[6997];
@(posedge clk);
#1;data_in = testData5[6998];
@(posedge clk);
#1;data_in = testData5[6999];
@(posedge clk);
#1;data_in = testData5[7000];
@(posedge clk);
#1;data_in = testData5[7001];
@(posedge clk);
#1;data_in = testData5[7002];
@(posedge clk);
#1;data_in = testData5[7003];
@(posedge clk);
#1;data_in = testData5[7004];
@(posedge clk);
#1;data_in = testData5[7005];
@(posedge clk);
#1;data_in = testData5[7006];
@(posedge clk);
#1;data_in = testData5[7007];
@(posedge clk);
#1;data_in = testData5[7008];
@(posedge clk);
#1;data_in = testData5[7009];
@(posedge clk);
#1;data_in = testData5[7010];
@(posedge clk);
#1;data_in = testData5[7011];
@(posedge clk);
#1;data_in = testData5[7012];
@(posedge clk);
#1;data_in = testData5[7013];
@(posedge clk);
#1;data_in = testData5[7014];
@(posedge clk);
#1;data_in = testData5[7015];
@(posedge clk);
#1;data_in = testData5[7016];
@(posedge clk);
#1;data_in = testData5[7017];
@(posedge clk);
#1;data_in = testData5[7018];
@(posedge clk);
#1;data_in = testData5[7019];
@(posedge clk);
#1;data_in = testData5[7020];
@(posedge clk);
#1;data_in = testData5[7021];
@(posedge clk);
#1;data_in = testData5[7022];
@(posedge clk);
#1;data_in = testData5[7023];
@(posedge clk);
#1;data_in = testData5[7024];
@(posedge clk);
#1;data_in = testData5[7025];
@(posedge clk);
#1;data_in = testData5[7026];
@(posedge clk);
#1;data_in = testData5[7027];
@(posedge clk);
#1;data_in = testData5[7028];
@(posedge clk);
#1;data_in = testData5[7029];
@(posedge clk);
#1;data_in = testData5[7030];
@(posedge clk);
#1;data_in = testData5[7031];
@(posedge clk);
#1;data_in = testData5[7032];
@(posedge clk);
#1;data_in = testData5[7033];
@(posedge clk);
#1;data_in = testData5[7034];
@(posedge clk);
#1;data_in = testData5[7035];
@(posedge clk);
#1;data_in = testData5[7036];
@(posedge clk);
#1;data_in = testData5[7037];
@(posedge clk);
#1;data_in = testData5[7038];
@(posedge clk);
#1;data_in = testData5[7039];
@(posedge clk);
#1;data_in = testData5[7040];
@(posedge clk);
#1;data_in = testData5[7041];
@(posedge clk);
#1;data_in = testData5[7042];
@(posedge clk);
#1;data_in = testData5[7043];
@(posedge clk);
#1;data_in = testData5[7044];
@(posedge clk);
#1;data_in = testData5[7045];
@(posedge clk);
#1;data_in = testData5[7046];
@(posedge clk);
#1;data_in = testData5[7047];
@(posedge clk);
#1;data_in = testData5[7048];
@(posedge clk);
#1;data_in = testData5[7049];
@(posedge clk);
#1;data_in = testData5[7050];
@(posedge clk);
#1;data_in = testData5[7051];
@(posedge clk);
#1;data_in = testData5[7052];
@(posedge clk);
#1;data_in = testData5[7053];
@(posedge clk);
#1;data_in = testData5[7054];
@(posedge clk);
#1;data_in = testData5[7055];
@(posedge clk);
#1;data_in = testData5[7056];
@(posedge clk);
#1;data_in = testData5[7057];
@(posedge clk);
#1;data_in = testData5[7058];
@(posedge clk);
#1;data_in = testData5[7059];
@(posedge clk);
#1;data_in = testData5[7060];
@(posedge clk);
#1;data_in = testData5[7061];
@(posedge clk);
#1;data_in = testData5[7062];
@(posedge clk);
#1;data_in = testData5[7063];
@(posedge clk);
#1;data_in = testData5[7064];
@(posedge clk);
#1;data_in = testData5[7065];
@(posedge clk);
#1;data_in = testData5[7066];
@(posedge clk);
#1;data_in = testData5[7067];
@(posedge clk);
#1;data_in = testData5[7068];
@(posedge clk);
#1;data_in = testData5[7069];
@(posedge clk);
#1;data_in = testData5[7070];
@(posedge clk);
#1;data_in = testData5[7071];
@(posedge clk);
#1;data_in = testData5[7072];
@(posedge clk);
#1;data_in = testData5[7073];
@(posedge clk);
#1;data_in = testData5[7074];
@(posedge clk);
#1;data_in = testData5[7075];
@(posedge clk);
#1;data_in = testData5[7076];
@(posedge clk);
#1;data_in = testData5[7077];
@(posedge clk);
#1;data_in = testData5[7078];
@(posedge clk);
#1;data_in = testData5[7079];
@(posedge clk);
#1;data_in = testData5[7080];
@(posedge clk);
#1;data_in = testData5[7081];
@(posedge clk);
#1;data_in = testData5[7082];
@(posedge clk);
#1;data_in = testData5[7083];
@(posedge clk);
#1;data_in = testData5[7084];
@(posedge clk);
#1;data_in = testData5[7085];
@(posedge clk);
#1;data_in = testData5[7086];
@(posedge clk);
#1;data_in = testData5[7087];
@(posedge clk);
#1;data_in = testData5[7088];
@(posedge clk);
#1;data_in = testData5[7089];
@(posedge clk);
#1;data_in = testData5[7090];
@(posedge clk);
#1;data_in = testData5[7091];
@(posedge clk);
#1;data_in = testData5[7092];
@(posedge clk);
#1;data_in = testData5[7093];
@(posedge clk);
#1;data_in = testData5[7094];
@(posedge clk);
#1;data_in = testData5[7095];
@(posedge clk);
#1;data_in = testData5[7096];
@(posedge clk);
#1;data_in = testData5[7097];
@(posedge clk);
#1;data_in = testData5[7098];
@(posedge clk);
#1;data_in = testData5[7099];
@(posedge clk);
#1;data_in = testData5[7100];
@(posedge clk);
#1;data_in = testData5[7101];
@(posedge clk);
#1;data_in = testData5[7102];
@(posedge clk);
#1;data_in = testData5[7103];
@(posedge clk);
#1;data_in = testData5[7104];
@(posedge clk);
#1;data_in = testData5[7105];
@(posedge clk);
#1;data_in = testData5[7106];
@(posedge clk);
#1;data_in = testData5[7107];
@(posedge clk);
#1;data_in = testData5[7108];
@(posedge clk);
#1;data_in = testData5[7109];
@(posedge clk);
#1;data_in = testData5[7110];
@(posedge clk);
#1;data_in = testData5[7111];
@(posedge clk);
#1;data_in = testData5[7112];
@(posedge clk);
#1;data_in = testData5[7113];
@(posedge clk);
#1;data_in = testData5[7114];
@(posedge clk);
#1;data_in = testData5[7115];
@(posedge clk);
#1;data_in = testData5[7116];
@(posedge clk);
#1;data_in = testData5[7117];
@(posedge clk);
#1;data_in = testData5[7118];
@(posedge clk);
#1;data_in = testData5[7119];
@(posedge clk);
#1;data_in = testData5[7120];
@(posedge clk);
#1;data_in = testData5[7121];
@(posedge clk);
#1;data_in = testData5[7122];
@(posedge clk);
#1;data_in = testData5[7123];
@(posedge clk);
#1;data_in = testData5[7124];
@(posedge clk);
#1;data_in = testData5[7125];
@(posedge clk);
#1;data_in = testData5[7126];
@(posedge clk);
#1;data_in = testData5[7127];
@(posedge clk);
#1;data_in = testData5[7128];
@(posedge clk);
#1;data_in = testData5[7129];
@(posedge clk);
#1;data_in = testData5[7130];
@(posedge clk);
#1;data_in = testData5[7131];
@(posedge clk);
#1;data_in = testData5[7132];
@(posedge clk);
#1;data_in = testData5[7133];
@(posedge clk);
#1;data_in = testData5[7134];
@(posedge clk);
#1;data_in = testData5[7135];
@(posedge clk);
#1;data_in = testData5[7136];
@(posedge clk);
#1;data_in = testData5[7137];
@(posedge clk);
#1;data_in = testData5[7138];
@(posedge clk);
#1;data_in = testData5[7139];
@(posedge clk);
#1;data_in = testData5[7140];
@(posedge clk);
#1;data_in = testData5[7141];
@(posedge clk);
#1;data_in = testData5[7142];
@(posedge clk);
#1;data_in = testData5[7143];
@(posedge clk);
#1;data_in = testData5[7144];
@(posedge clk);
#1;data_in = testData5[7145];
@(posedge clk);
#1;data_in = testData5[7146];
@(posedge clk);
#1;data_in = testData5[7147];
@(posedge clk);
#1;data_in = testData5[7148];
@(posedge clk);
#1;data_in = testData5[7149];
@(posedge clk);
#1;data_in = testData5[7150];
@(posedge clk);
#1;data_in = testData5[7151];
@(posedge clk);
#1;data_in = testData5[7152];
@(posedge clk);
#1;data_in = testData5[7153];
@(posedge clk);
#1;data_in = testData5[7154];
@(posedge clk);
#1;data_in = testData5[7155];
@(posedge clk);
#1;data_in = testData5[7156];
@(posedge clk);
#1;data_in = testData5[7157];
@(posedge clk);
#1;data_in = testData5[7158];
@(posedge clk);
#1;data_in = testData5[7159];
@(posedge clk);
#1;data_in = testData5[7160];
@(posedge clk);
#1;data_in = testData5[7161];
@(posedge clk);
#1;data_in = testData5[7162];
@(posedge clk);
#1;data_in = testData5[7163];
@(posedge clk);
#1;data_in = testData5[7164];
@(posedge clk);
#1;data_in = testData5[7165];
@(posedge clk);
#1;data_in = testData5[7166];
@(posedge clk);
#1;data_in = testData5[7167];
@(posedge clk);
#1;data_in = testData5[7168];
@(posedge clk);
#1;data_in = testData5[7169];
@(posedge clk);
#1;data_in = testData5[7170];
@(posedge clk);
#1;data_in = testData5[7171];
@(posedge clk);
#1;data_in = testData5[7172];
@(posedge clk);
#1;data_in = testData5[7173];
@(posedge clk);
#1;data_in = testData5[7174];
@(posedge clk);
#1;data_in = testData5[7175];
@(posedge clk);
#1;data_in = testData5[7176];
@(posedge clk);
#1;data_in = testData5[7177];
@(posedge clk);
#1;data_in = testData5[7178];
@(posedge clk);
#1;data_in = testData5[7179];
@(posedge clk);
#1;data_in = testData5[7180];
@(posedge clk);
#1;data_in = testData5[7181];
@(posedge clk);
#1;data_in = testData5[7182];
@(posedge clk);
#1;data_in = testData5[7183];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[7184]; 
@(posedge clk);
#1;data_in = testData5[7185];
@(posedge clk);
#1;data_in = testData5[7186];
@(posedge clk);
#1;data_in = testData5[7187];
@(posedge clk);
#1;data_in = testData5[7188];
@(posedge clk);
#1;data_in = testData5[7189];
@(posedge clk);
#1;data_in = testData5[7190];
@(posedge clk);
#1;data_in = testData5[7191];
@(posedge clk);
#1;data_in = testData5[7192];
@(posedge clk);
#1;data_in = testData5[7193];
@(posedge clk);
#1;data_in = testData5[7194];
@(posedge clk);
#1;data_in = testData5[7195];
@(posedge clk);
#1;data_in = testData5[7196];
@(posedge clk);
#1;data_in = testData5[7197];
@(posedge clk);
#1;data_in = testData5[7198];
@(posedge clk);
#1;data_in = testData5[7199];
@(posedge clk);
#1;data_in = testData5[7200];
@(posedge clk);
#1;data_in = testData5[7201];
@(posedge clk);
#1;data_in = testData5[7202];
@(posedge clk);
#1;data_in = testData5[7203];
@(posedge clk);
#1;data_in = testData5[7204];
@(posedge clk);
#1;data_in = testData5[7205];
@(posedge clk);
#1;data_in = testData5[7206];
@(posedge clk);
#1;data_in = testData5[7207];
@(posedge clk);
#1;data_in = testData5[7208];
@(posedge clk);
#1;data_in = testData5[7209];
@(posedge clk);
#1;data_in = testData5[7210];
@(posedge clk);
#1;data_in = testData5[7211];
@(posedge clk);
#1;data_in = testData5[7212];
@(posedge clk);
#1;data_in = testData5[7213];
@(posedge clk);
#1;data_in = testData5[7214];
@(posedge clk);
#1;data_in = testData5[7215];
@(posedge clk);
#1;data_in = testData5[7216];
@(posedge clk);
#1;data_in = testData5[7217];
@(posedge clk);
#1;data_in = testData5[7218];
@(posedge clk);
#1;data_in = testData5[7219];
@(posedge clk);
#1;data_in = testData5[7220];
@(posedge clk);
#1;data_in = testData5[7221];
@(posedge clk);
#1;data_in = testData5[7222];
@(posedge clk);
#1;data_in = testData5[7223];
@(posedge clk);
#1;data_in = testData5[7224];
@(posedge clk);
#1;data_in = testData5[7225];
@(posedge clk);
#1;data_in = testData5[7226];
@(posedge clk);
#1;data_in = testData5[7227];
@(posedge clk);
#1;data_in = testData5[7228];
@(posedge clk);
#1;data_in = testData5[7229];
@(posedge clk);
#1;data_in = testData5[7230];
@(posedge clk);
#1;data_in = testData5[7231];
@(posedge clk);
#1;data_in = testData5[7232];
@(posedge clk);
#1;data_in = testData5[7233];
@(posedge clk);
#1;data_in = testData5[7234];
@(posedge clk);
#1;data_in = testData5[7235];
@(posedge clk);
#1;data_in = testData5[7236];
@(posedge clk);
#1;data_in = testData5[7237];
@(posedge clk);
#1;data_in = testData5[7238];
@(posedge clk);
#1;data_in = testData5[7239];
@(posedge clk);
#1;data_in = testData5[7240];
@(posedge clk);
#1;data_in = testData5[7241];
@(posedge clk);
#1;data_in = testData5[7242];
@(posedge clk);
#1;data_in = testData5[7243];
@(posedge clk);
#1;data_in = testData5[7244];
@(posedge clk);
#1;data_in = testData5[7245];
@(posedge clk);
#1;data_in = testData5[7246];
@(posedge clk);
#1;data_in = testData5[7247];
@(posedge clk);
#1;data_in = testData5[7248];
@(posedge clk);
#1;data_in = testData5[7249];
@(posedge clk);
#1;data_in = testData5[7250];
@(posedge clk);
#1;data_in = testData5[7251];
@(posedge clk);
#1;data_in = testData5[7252];
@(posedge clk);
#1;data_in = testData5[7253];
@(posedge clk);
#1;data_in = testData5[7254];
@(posedge clk);
#1;data_in = testData5[7255];
@(posedge clk);
#1;data_in = testData5[7256];
@(posedge clk);
#1;data_in = testData5[7257];
@(posedge clk);
#1;data_in = testData5[7258];
@(posedge clk);
#1;data_in = testData5[7259];
@(posedge clk);
#1;data_in = testData5[7260];
@(posedge clk);
#1;data_in = testData5[7261];
@(posedge clk);
#1;data_in = testData5[7262];
@(posedge clk);
#1;data_in = testData5[7263];
@(posedge clk);
#1;data_in = testData5[7264];
@(posedge clk);
#1;data_in = testData5[7265];
@(posedge clk);
#1;data_in = testData5[7266];
@(posedge clk);
#1;data_in = testData5[7267];
@(posedge clk);
#1;data_in = testData5[7268];
@(posedge clk);
#1;data_in = testData5[7269];
@(posedge clk);
#1;data_in = testData5[7270];
@(posedge clk);
#1;data_in = testData5[7271];
@(posedge clk);
#1;data_in = testData5[7272];
@(posedge clk);
#1;data_in = testData5[7273];
@(posedge clk);
#1;data_in = testData5[7274];
@(posedge clk);
#1;data_in = testData5[7275];
@(posedge clk);
#1;data_in = testData5[7276];
@(posedge clk);
#1;data_in = testData5[7277];
@(posedge clk);
#1;data_in = testData5[7278];
@(posedge clk);
#1;data_in = testData5[7279];
@(posedge clk);
#1;data_in = testData5[7280];
@(posedge clk);
#1;data_in = testData5[7281];
@(posedge clk);
#1;data_in = testData5[7282];
@(posedge clk);
#1;data_in = testData5[7283];
@(posedge clk);
#1;data_in = testData5[7284];
@(posedge clk);
#1;data_in = testData5[7285];
@(posedge clk);
#1;data_in = testData5[7286];
@(posedge clk);
#1;data_in = testData5[7287];
@(posedge clk);
#1;data_in = testData5[7288];
@(posedge clk);
#1;data_in = testData5[7289];
@(posedge clk);
#1;data_in = testData5[7290];
@(posedge clk);
#1;data_in = testData5[7291];
@(posedge clk);
#1;data_in = testData5[7292];
@(posedge clk);
#1;data_in = testData5[7293];
@(posedge clk);
#1;data_in = testData5[7294];
@(posedge clk);
#1;data_in = testData5[7295];
@(posedge clk);
#1;data_in = testData5[7296];
@(posedge clk);
#1;data_in = testData5[7297];
@(posedge clk);
#1;data_in = testData5[7298];
@(posedge clk);
#1;data_in = testData5[7299];
@(posedge clk);
#1;data_in = testData5[7300];
@(posedge clk);
#1;data_in = testData5[7301];
@(posedge clk);
#1;data_in = testData5[7302];
@(posedge clk);
#1;data_in = testData5[7303];
@(posedge clk);
#1;data_in = testData5[7304];
@(posedge clk);
#1;data_in = testData5[7305];
@(posedge clk);
#1;data_in = testData5[7306];
@(posedge clk);
#1;data_in = testData5[7307];
@(posedge clk);
#1;data_in = testData5[7308];
@(posedge clk);
#1;data_in = testData5[7309];
@(posedge clk);
#1;data_in = testData5[7310];
@(posedge clk);
#1;data_in = testData5[7311];
@(posedge clk);
#1;data_in = testData5[7312];
@(posedge clk);
#1;data_in = testData5[7313];
@(posedge clk);
#1;data_in = testData5[7314];
@(posedge clk);
#1;data_in = testData5[7315];
@(posedge clk);
#1;data_in = testData5[7316];
@(posedge clk);
#1;data_in = testData5[7317];
@(posedge clk);
#1;data_in = testData5[7318];
@(posedge clk);
#1;data_in = testData5[7319];
@(posedge clk);
#1;data_in = testData5[7320];
@(posedge clk);
#1;data_in = testData5[7321];
@(posedge clk);
#1;data_in = testData5[7322];
@(posedge clk);
#1;data_in = testData5[7323];
@(posedge clk);
#1;data_in = testData5[7324];
@(posedge clk);
#1;data_in = testData5[7325];
@(posedge clk);
#1;data_in = testData5[7326];
@(posedge clk);
#1;data_in = testData5[7327];
@(posedge clk);
#1;data_in = testData5[7328];
@(posedge clk);
#1;data_in = testData5[7329];
@(posedge clk);
#1;data_in = testData5[7330];
@(posedge clk);
#1;data_in = testData5[7331];
@(posedge clk);
#1;data_in = testData5[7332];
@(posedge clk);
#1;data_in = testData5[7333];
@(posedge clk);
#1;data_in = testData5[7334];
@(posedge clk);
#1;data_in = testData5[7335];
@(posedge clk);
#1;data_in = testData5[7336];
@(posedge clk);
#1;data_in = testData5[7337];
@(posedge clk);
#1;data_in = testData5[7338];
@(posedge clk);
#1;data_in = testData5[7339];
@(posedge clk);
#1;data_in = testData5[7340];
@(posedge clk);
#1;data_in = testData5[7341];
@(posedge clk);
#1;data_in = testData5[7342];
@(posedge clk);
#1;data_in = testData5[7343];
@(posedge clk);
#1;data_in = testData5[7344];
@(posedge clk);
#1;data_in = testData5[7345];
@(posedge clk);
#1;data_in = testData5[7346];
@(posedge clk);
#1;data_in = testData5[7347];
@(posedge clk);
#1;data_in = testData5[7348];
@(posedge clk);
#1;data_in = testData5[7349];
@(posedge clk);
#1;data_in = testData5[7350];
@(posedge clk);
#1;data_in = testData5[7351];
@(posedge clk);
#1;data_in = testData5[7352];
@(posedge clk);
#1;data_in = testData5[7353];
@(posedge clk);
#1;data_in = testData5[7354];
@(posedge clk);
#1;data_in = testData5[7355];
@(posedge clk);
#1;data_in = testData5[7356];
@(posedge clk);
#1;data_in = testData5[7357];
@(posedge clk);
#1;data_in = testData5[7358];
@(posedge clk);
#1;data_in = testData5[7359];
@(posedge clk);
#1;data_in = testData5[7360];
@(posedge clk);
#1;data_in = testData5[7361];
@(posedge clk);
#1;data_in = testData5[7362];
@(posedge clk);
#1;data_in = testData5[7363];
@(posedge clk);
#1;data_in = testData5[7364];
@(posedge clk);
#1;data_in = testData5[7365];
@(posedge clk);
#1;data_in = testData5[7366];
@(posedge clk);
#1;data_in = testData5[7367];
@(posedge clk);
#1;data_in = testData5[7368];
@(posedge clk);
#1;data_in = testData5[7369];
@(posedge clk);
#1;data_in = testData5[7370];
@(posedge clk);
#1;data_in = testData5[7371];
@(posedge clk);
#1;data_in = testData5[7372];
@(posedge clk);
#1;data_in = testData5[7373];
@(posedge clk);
#1;data_in = testData5[7374];
@(posedge clk);
#1;data_in = testData5[7375];
@(posedge clk);
#1;data_in = testData5[7376];
@(posedge clk);
#1;data_in = testData5[7377];
@(posedge clk);
#1;data_in = testData5[7378];
@(posedge clk);
#1;data_in = testData5[7379];
@(posedge clk);
#1;data_in = testData5[7380];
@(posedge clk);
#1;data_in = testData5[7381];
@(posedge clk);
#1;data_in = testData5[7382];
@(posedge clk);
#1;data_in = testData5[7383];
@(posedge clk);
#1;data_in = testData5[7384];
@(posedge clk);
#1;data_in = testData5[7385];
@(posedge clk);
#1;data_in = testData5[7386];
@(posedge clk);
#1;data_in = testData5[7387];
@(posedge clk);
#1;data_in = testData5[7388];
@(posedge clk);
#1;data_in = testData5[7389];
@(posedge clk);
#1;data_in = testData5[7390];
@(posedge clk);
#1;data_in = testData5[7391];
@(posedge clk);
#1;data_in = testData5[7392];
@(posedge clk);
#1;data_in = testData5[7393];
@(posedge clk);
#1;data_in = testData5[7394];
@(posedge clk);
#1;data_in = testData5[7395];
@(posedge clk);
#1;data_in = testData5[7396];
@(posedge clk);
#1;data_in = testData5[7397];
@(posedge clk);
#1;data_in = testData5[7398];
@(posedge clk);
#1;data_in = testData5[7399];
@(posedge clk);
#1;data_in = testData5[7400];
@(posedge clk);
#1;data_in = testData5[7401];
@(posedge clk);
#1;data_in = testData5[7402];
@(posedge clk);
#1;data_in = testData5[7403];
@(posedge clk);
#1;data_in = testData5[7404];
@(posedge clk);
#1;data_in = testData5[7405];
@(posedge clk);
#1;data_in = testData5[7406];
@(posedge clk);
#1;data_in = testData5[7407];
@(posedge clk);
#1;data_in = testData5[7408];
@(posedge clk);
#1;data_in = testData5[7409];
@(posedge clk);
#1;data_in = testData5[7410];
@(posedge clk);
#1;data_in = testData5[7411];
@(posedge clk);
#1;data_in = testData5[7412];
@(posedge clk);
#1;data_in = testData5[7413];
@(posedge clk);
#1;data_in = testData5[7414];
@(posedge clk);
#1;data_in = testData5[7415];
@(posedge clk);
#1;data_in = testData5[7416];
@(posedge clk);
#1;data_in = testData5[7417];
@(posedge clk);
#1;data_in = testData5[7418];
@(posedge clk);
#1;data_in = testData5[7419];
@(posedge clk);
#1;data_in = testData5[7420];
@(posedge clk);
#1;data_in = testData5[7421];
@(posedge clk);
#1;data_in = testData5[7422];
@(posedge clk);
#1;data_in = testData5[7423];
@(posedge clk);
#1;data_in = testData5[7424];
@(posedge clk);
#1;data_in = testData5[7425];
@(posedge clk);
#1;data_in = testData5[7426];
@(posedge clk);
#1;data_in = testData5[7427];
@(posedge clk);
#1;data_in = testData5[7428];
@(posedge clk);
#1;data_in = testData5[7429];
@(posedge clk);
#1;data_in = testData5[7430];
@(posedge clk);
#1;data_in = testData5[7431];
@(posedge clk);
#1;data_in = testData5[7432];
@(posedge clk);
#1;data_in = testData5[7433];
@(posedge clk);
#1;data_in = testData5[7434];
@(posedge clk);
#1;data_in = testData5[7435];
@(posedge clk);
#1;data_in = testData5[7436];
@(posedge clk);
#1;data_in = testData5[7437];
@(posedge clk);
#1;data_in = testData5[7438];
@(posedge clk);
#1;data_in = testData5[7439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[7440]; 
@(posedge clk);
#1;data_in = testData5[7441];
@(posedge clk);
#1;data_in = testData5[7442];
@(posedge clk);
#1;data_in = testData5[7443];
@(posedge clk);
#1;data_in = testData5[7444];
@(posedge clk);
#1;data_in = testData5[7445];
@(posedge clk);
#1;data_in = testData5[7446];
@(posedge clk);
#1;data_in = testData5[7447];
@(posedge clk);
#1;data_in = testData5[7448];
@(posedge clk);
#1;data_in = testData5[7449];
@(posedge clk);
#1;data_in = testData5[7450];
@(posedge clk);
#1;data_in = testData5[7451];
@(posedge clk);
#1;data_in = testData5[7452];
@(posedge clk);
#1;data_in = testData5[7453];
@(posedge clk);
#1;data_in = testData5[7454];
@(posedge clk);
#1;data_in = testData5[7455];
@(posedge clk);
#1;data_in = testData5[7456];
@(posedge clk);
#1;data_in = testData5[7457];
@(posedge clk);
#1;data_in = testData5[7458];
@(posedge clk);
#1;data_in = testData5[7459];
@(posedge clk);
#1;data_in = testData5[7460];
@(posedge clk);
#1;data_in = testData5[7461];
@(posedge clk);
#1;data_in = testData5[7462];
@(posedge clk);
#1;data_in = testData5[7463];
@(posedge clk);
#1;data_in = testData5[7464];
@(posedge clk);
#1;data_in = testData5[7465];
@(posedge clk);
#1;data_in = testData5[7466];
@(posedge clk);
#1;data_in = testData5[7467];
@(posedge clk);
#1;data_in = testData5[7468];
@(posedge clk);
#1;data_in = testData5[7469];
@(posedge clk);
#1;data_in = testData5[7470];
@(posedge clk);
#1;data_in = testData5[7471];
@(posedge clk);
#1;data_in = testData5[7472];
@(posedge clk);
#1;data_in = testData5[7473];
@(posedge clk);
#1;data_in = testData5[7474];
@(posedge clk);
#1;data_in = testData5[7475];
@(posedge clk);
#1;data_in = testData5[7476];
@(posedge clk);
#1;data_in = testData5[7477];
@(posedge clk);
#1;data_in = testData5[7478];
@(posedge clk);
#1;data_in = testData5[7479];
@(posedge clk);
#1;data_in = testData5[7480];
@(posedge clk);
#1;data_in = testData5[7481];
@(posedge clk);
#1;data_in = testData5[7482];
@(posedge clk);
#1;data_in = testData5[7483];
@(posedge clk);
#1;data_in = testData5[7484];
@(posedge clk);
#1;data_in = testData5[7485];
@(posedge clk);
#1;data_in = testData5[7486];
@(posedge clk);
#1;data_in = testData5[7487];
@(posedge clk);
#1;data_in = testData5[7488];
@(posedge clk);
#1;data_in = testData5[7489];
@(posedge clk);
#1;data_in = testData5[7490];
@(posedge clk);
#1;data_in = testData5[7491];
@(posedge clk);
#1;data_in = testData5[7492];
@(posedge clk);
#1;data_in = testData5[7493];
@(posedge clk);
#1;data_in = testData5[7494];
@(posedge clk);
#1;data_in = testData5[7495];
@(posedge clk);
#1;data_in = testData5[7496];
@(posedge clk);
#1;data_in = testData5[7497];
@(posedge clk);
#1;data_in = testData5[7498];
@(posedge clk);
#1;data_in = testData5[7499];
@(posedge clk);
#1;data_in = testData5[7500];
@(posedge clk);
#1;data_in = testData5[7501];
@(posedge clk);
#1;data_in = testData5[7502];
@(posedge clk);
#1;data_in = testData5[7503];
@(posedge clk);
#1;data_in = testData5[7504];
@(posedge clk);
#1;data_in = testData5[7505];
@(posedge clk);
#1;data_in = testData5[7506];
@(posedge clk);
#1;data_in = testData5[7507];
@(posedge clk);
#1;data_in = testData5[7508];
@(posedge clk);
#1;data_in = testData5[7509];
@(posedge clk);
#1;data_in = testData5[7510];
@(posedge clk);
#1;data_in = testData5[7511];
@(posedge clk);
#1;data_in = testData5[7512];
@(posedge clk);
#1;data_in = testData5[7513];
@(posedge clk);
#1;data_in = testData5[7514];
@(posedge clk);
#1;data_in = testData5[7515];
@(posedge clk);
#1;data_in = testData5[7516];
@(posedge clk);
#1;data_in = testData5[7517];
@(posedge clk);
#1;data_in = testData5[7518];
@(posedge clk);
#1;data_in = testData5[7519];
@(posedge clk);
#1;data_in = testData5[7520];
@(posedge clk);
#1;data_in = testData5[7521];
@(posedge clk);
#1;data_in = testData5[7522];
@(posedge clk);
#1;data_in = testData5[7523];
@(posedge clk);
#1;data_in = testData5[7524];
@(posedge clk);
#1;data_in = testData5[7525];
@(posedge clk);
#1;data_in = testData5[7526];
@(posedge clk);
#1;data_in = testData5[7527];
@(posedge clk);
#1;data_in = testData5[7528];
@(posedge clk);
#1;data_in = testData5[7529];
@(posedge clk);
#1;data_in = testData5[7530];
@(posedge clk);
#1;data_in = testData5[7531];
@(posedge clk);
#1;data_in = testData5[7532];
@(posedge clk);
#1;data_in = testData5[7533];
@(posedge clk);
#1;data_in = testData5[7534];
@(posedge clk);
#1;data_in = testData5[7535];
@(posedge clk);
#1;data_in = testData5[7536];
@(posedge clk);
#1;data_in = testData5[7537];
@(posedge clk);
#1;data_in = testData5[7538];
@(posedge clk);
#1;data_in = testData5[7539];
@(posedge clk);
#1;data_in = testData5[7540];
@(posedge clk);
#1;data_in = testData5[7541];
@(posedge clk);
#1;data_in = testData5[7542];
@(posedge clk);
#1;data_in = testData5[7543];
@(posedge clk);
#1;data_in = testData5[7544];
@(posedge clk);
#1;data_in = testData5[7545];
@(posedge clk);
#1;data_in = testData5[7546];
@(posedge clk);
#1;data_in = testData5[7547];
@(posedge clk);
#1;data_in = testData5[7548];
@(posedge clk);
#1;data_in = testData5[7549];
@(posedge clk);
#1;data_in = testData5[7550];
@(posedge clk);
#1;data_in = testData5[7551];
@(posedge clk);
#1;data_in = testData5[7552];
@(posedge clk);
#1;data_in = testData5[7553];
@(posedge clk);
#1;data_in = testData5[7554];
@(posedge clk);
#1;data_in = testData5[7555];
@(posedge clk);
#1;data_in = testData5[7556];
@(posedge clk);
#1;data_in = testData5[7557];
@(posedge clk);
#1;data_in = testData5[7558];
@(posedge clk);
#1;data_in = testData5[7559];
@(posedge clk);
#1;data_in = testData5[7560];
@(posedge clk);
#1;data_in = testData5[7561];
@(posedge clk);
#1;data_in = testData5[7562];
@(posedge clk);
#1;data_in = testData5[7563];
@(posedge clk);
#1;data_in = testData5[7564];
@(posedge clk);
#1;data_in = testData5[7565];
@(posedge clk);
#1;data_in = testData5[7566];
@(posedge clk);
#1;data_in = testData5[7567];
@(posedge clk);
#1;data_in = testData5[7568];
@(posedge clk);
#1;data_in = testData5[7569];
@(posedge clk);
#1;data_in = testData5[7570];
@(posedge clk);
#1;data_in = testData5[7571];
@(posedge clk);
#1;data_in = testData5[7572];
@(posedge clk);
#1;data_in = testData5[7573];
@(posedge clk);
#1;data_in = testData5[7574];
@(posedge clk);
#1;data_in = testData5[7575];
@(posedge clk);
#1;data_in = testData5[7576];
@(posedge clk);
#1;data_in = testData5[7577];
@(posedge clk);
#1;data_in = testData5[7578];
@(posedge clk);
#1;data_in = testData5[7579];
@(posedge clk);
#1;data_in = testData5[7580];
@(posedge clk);
#1;data_in = testData5[7581];
@(posedge clk);
#1;data_in = testData5[7582];
@(posedge clk);
#1;data_in = testData5[7583];
@(posedge clk);
#1;data_in = testData5[7584];
@(posedge clk);
#1;data_in = testData5[7585];
@(posedge clk);
#1;data_in = testData5[7586];
@(posedge clk);
#1;data_in = testData5[7587];
@(posedge clk);
#1;data_in = testData5[7588];
@(posedge clk);
#1;data_in = testData5[7589];
@(posedge clk);
#1;data_in = testData5[7590];
@(posedge clk);
#1;data_in = testData5[7591];
@(posedge clk);
#1;data_in = testData5[7592];
@(posedge clk);
#1;data_in = testData5[7593];
@(posedge clk);
#1;data_in = testData5[7594];
@(posedge clk);
#1;data_in = testData5[7595];
@(posedge clk);
#1;data_in = testData5[7596];
@(posedge clk);
#1;data_in = testData5[7597];
@(posedge clk);
#1;data_in = testData5[7598];
@(posedge clk);
#1;data_in = testData5[7599];
@(posedge clk);
#1;data_in = testData5[7600];
@(posedge clk);
#1;data_in = testData5[7601];
@(posedge clk);
#1;data_in = testData5[7602];
@(posedge clk);
#1;data_in = testData5[7603];
@(posedge clk);
#1;data_in = testData5[7604];
@(posedge clk);
#1;data_in = testData5[7605];
@(posedge clk);
#1;data_in = testData5[7606];
@(posedge clk);
#1;data_in = testData5[7607];
@(posedge clk);
#1;data_in = testData5[7608];
@(posedge clk);
#1;data_in = testData5[7609];
@(posedge clk);
#1;data_in = testData5[7610];
@(posedge clk);
#1;data_in = testData5[7611];
@(posedge clk);
#1;data_in = testData5[7612];
@(posedge clk);
#1;data_in = testData5[7613];
@(posedge clk);
#1;data_in = testData5[7614];
@(posedge clk);
#1;data_in = testData5[7615];
@(posedge clk);
#1;data_in = testData5[7616];
@(posedge clk);
#1;data_in = testData5[7617];
@(posedge clk);
#1;data_in = testData5[7618];
@(posedge clk);
#1;data_in = testData5[7619];
@(posedge clk);
#1;data_in = testData5[7620];
@(posedge clk);
#1;data_in = testData5[7621];
@(posedge clk);
#1;data_in = testData5[7622];
@(posedge clk);
#1;data_in = testData5[7623];
@(posedge clk);
#1;data_in = testData5[7624];
@(posedge clk);
#1;data_in = testData5[7625];
@(posedge clk);
#1;data_in = testData5[7626];
@(posedge clk);
#1;data_in = testData5[7627];
@(posedge clk);
#1;data_in = testData5[7628];
@(posedge clk);
#1;data_in = testData5[7629];
@(posedge clk);
#1;data_in = testData5[7630];
@(posedge clk);
#1;data_in = testData5[7631];
@(posedge clk);
#1;data_in = testData5[7632];
@(posedge clk);
#1;data_in = testData5[7633];
@(posedge clk);
#1;data_in = testData5[7634];
@(posedge clk);
#1;data_in = testData5[7635];
@(posedge clk);
#1;data_in = testData5[7636];
@(posedge clk);
#1;data_in = testData5[7637];
@(posedge clk);
#1;data_in = testData5[7638];
@(posedge clk);
#1;data_in = testData5[7639];
@(posedge clk);
#1;data_in = testData5[7640];
@(posedge clk);
#1;data_in = testData5[7641];
@(posedge clk);
#1;data_in = testData5[7642];
@(posedge clk);
#1;data_in = testData5[7643];
@(posedge clk);
#1;data_in = testData5[7644];
@(posedge clk);
#1;data_in = testData5[7645];
@(posedge clk);
#1;data_in = testData5[7646];
@(posedge clk);
#1;data_in = testData5[7647];
@(posedge clk);
#1;data_in = testData5[7648];
@(posedge clk);
#1;data_in = testData5[7649];
@(posedge clk);
#1;data_in = testData5[7650];
@(posedge clk);
#1;data_in = testData5[7651];
@(posedge clk);
#1;data_in = testData5[7652];
@(posedge clk);
#1;data_in = testData5[7653];
@(posedge clk);
#1;data_in = testData5[7654];
@(posedge clk);
#1;data_in = testData5[7655];
@(posedge clk);
#1;data_in = testData5[7656];
@(posedge clk);
#1;data_in = testData5[7657];
@(posedge clk);
#1;data_in = testData5[7658];
@(posedge clk);
#1;data_in = testData5[7659];
@(posedge clk);
#1;data_in = testData5[7660];
@(posedge clk);
#1;data_in = testData5[7661];
@(posedge clk);
#1;data_in = testData5[7662];
@(posedge clk);
#1;data_in = testData5[7663];
@(posedge clk);
#1;data_in = testData5[7664];
@(posedge clk);
#1;data_in = testData5[7665];
@(posedge clk);
#1;data_in = testData5[7666];
@(posedge clk);
#1;data_in = testData5[7667];
@(posedge clk);
#1;data_in = testData5[7668];
@(posedge clk);
#1;data_in = testData5[7669];
@(posedge clk);
#1;data_in = testData5[7670];
@(posedge clk);
#1;data_in = testData5[7671];
@(posedge clk);
#1;data_in = testData5[7672];
@(posedge clk);
#1;data_in = testData5[7673];
@(posedge clk);
#1;data_in = testData5[7674];
@(posedge clk);
#1;data_in = testData5[7675];
@(posedge clk);
#1;data_in = testData5[7676];
@(posedge clk);
#1;data_in = testData5[7677];
@(posedge clk);
#1;data_in = testData5[7678];
@(posedge clk);
#1;data_in = testData5[7679];
@(posedge clk);
#1;data_in = testData5[7680];
@(posedge clk);
#1;data_in = testData5[7681];
@(posedge clk);
#1;data_in = testData5[7682];
@(posedge clk);
#1;data_in = testData5[7683];
@(posedge clk);
#1;data_in = testData5[7684];
@(posedge clk);
#1;data_in = testData5[7685];
@(posedge clk);
#1;data_in = testData5[7686];
@(posedge clk);
#1;data_in = testData5[7687];
@(posedge clk);
#1;data_in = testData5[7688];
@(posedge clk);
#1;data_in = testData5[7689];
@(posedge clk);
#1;data_in = testData5[7690];
@(posedge clk);
#1;data_in = testData5[7691];
@(posedge clk);
#1;data_in = testData5[7692];
@(posedge clk);
#1;data_in = testData5[7693];
@(posedge clk);
#1;data_in = testData5[7694];
@(posedge clk);
#1;data_in = testData5[7695];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[7696]; 
@(posedge clk);
#1;data_in = testData5[7697];
@(posedge clk);
#1;data_in = testData5[7698];
@(posedge clk);
#1;data_in = testData5[7699];
@(posedge clk);
#1;data_in = testData5[7700];
@(posedge clk);
#1;data_in = testData5[7701];
@(posedge clk);
#1;data_in = testData5[7702];
@(posedge clk);
#1;data_in = testData5[7703];
@(posedge clk);
#1;data_in = testData5[7704];
@(posedge clk);
#1;data_in = testData5[7705];
@(posedge clk);
#1;data_in = testData5[7706];
@(posedge clk);
#1;data_in = testData5[7707];
@(posedge clk);
#1;data_in = testData5[7708];
@(posedge clk);
#1;data_in = testData5[7709];
@(posedge clk);
#1;data_in = testData5[7710];
@(posedge clk);
#1;data_in = testData5[7711];
@(posedge clk);
#1;data_in = testData5[7712];
@(posedge clk);
#1;data_in = testData5[7713];
@(posedge clk);
#1;data_in = testData5[7714];
@(posedge clk);
#1;data_in = testData5[7715];
@(posedge clk);
#1;data_in = testData5[7716];
@(posedge clk);
#1;data_in = testData5[7717];
@(posedge clk);
#1;data_in = testData5[7718];
@(posedge clk);
#1;data_in = testData5[7719];
@(posedge clk);
#1;data_in = testData5[7720];
@(posedge clk);
#1;data_in = testData5[7721];
@(posedge clk);
#1;data_in = testData5[7722];
@(posedge clk);
#1;data_in = testData5[7723];
@(posedge clk);
#1;data_in = testData5[7724];
@(posedge clk);
#1;data_in = testData5[7725];
@(posedge clk);
#1;data_in = testData5[7726];
@(posedge clk);
#1;data_in = testData5[7727];
@(posedge clk);
#1;data_in = testData5[7728];
@(posedge clk);
#1;data_in = testData5[7729];
@(posedge clk);
#1;data_in = testData5[7730];
@(posedge clk);
#1;data_in = testData5[7731];
@(posedge clk);
#1;data_in = testData5[7732];
@(posedge clk);
#1;data_in = testData5[7733];
@(posedge clk);
#1;data_in = testData5[7734];
@(posedge clk);
#1;data_in = testData5[7735];
@(posedge clk);
#1;data_in = testData5[7736];
@(posedge clk);
#1;data_in = testData5[7737];
@(posedge clk);
#1;data_in = testData5[7738];
@(posedge clk);
#1;data_in = testData5[7739];
@(posedge clk);
#1;data_in = testData5[7740];
@(posedge clk);
#1;data_in = testData5[7741];
@(posedge clk);
#1;data_in = testData5[7742];
@(posedge clk);
#1;data_in = testData5[7743];
@(posedge clk);
#1;data_in = testData5[7744];
@(posedge clk);
#1;data_in = testData5[7745];
@(posedge clk);
#1;data_in = testData5[7746];
@(posedge clk);
#1;data_in = testData5[7747];
@(posedge clk);
#1;data_in = testData5[7748];
@(posedge clk);
#1;data_in = testData5[7749];
@(posedge clk);
#1;data_in = testData5[7750];
@(posedge clk);
#1;data_in = testData5[7751];
@(posedge clk);
#1;data_in = testData5[7752];
@(posedge clk);
#1;data_in = testData5[7753];
@(posedge clk);
#1;data_in = testData5[7754];
@(posedge clk);
#1;data_in = testData5[7755];
@(posedge clk);
#1;data_in = testData5[7756];
@(posedge clk);
#1;data_in = testData5[7757];
@(posedge clk);
#1;data_in = testData5[7758];
@(posedge clk);
#1;data_in = testData5[7759];
@(posedge clk);
#1;data_in = testData5[7760];
@(posedge clk);
#1;data_in = testData5[7761];
@(posedge clk);
#1;data_in = testData5[7762];
@(posedge clk);
#1;data_in = testData5[7763];
@(posedge clk);
#1;data_in = testData5[7764];
@(posedge clk);
#1;data_in = testData5[7765];
@(posedge clk);
#1;data_in = testData5[7766];
@(posedge clk);
#1;data_in = testData5[7767];
@(posedge clk);
#1;data_in = testData5[7768];
@(posedge clk);
#1;data_in = testData5[7769];
@(posedge clk);
#1;data_in = testData5[7770];
@(posedge clk);
#1;data_in = testData5[7771];
@(posedge clk);
#1;data_in = testData5[7772];
@(posedge clk);
#1;data_in = testData5[7773];
@(posedge clk);
#1;data_in = testData5[7774];
@(posedge clk);
#1;data_in = testData5[7775];
@(posedge clk);
#1;data_in = testData5[7776];
@(posedge clk);
#1;data_in = testData5[7777];
@(posedge clk);
#1;data_in = testData5[7778];
@(posedge clk);
#1;data_in = testData5[7779];
@(posedge clk);
#1;data_in = testData5[7780];
@(posedge clk);
#1;data_in = testData5[7781];
@(posedge clk);
#1;data_in = testData5[7782];
@(posedge clk);
#1;data_in = testData5[7783];
@(posedge clk);
#1;data_in = testData5[7784];
@(posedge clk);
#1;data_in = testData5[7785];
@(posedge clk);
#1;data_in = testData5[7786];
@(posedge clk);
#1;data_in = testData5[7787];
@(posedge clk);
#1;data_in = testData5[7788];
@(posedge clk);
#1;data_in = testData5[7789];
@(posedge clk);
#1;data_in = testData5[7790];
@(posedge clk);
#1;data_in = testData5[7791];
@(posedge clk);
#1;data_in = testData5[7792];
@(posedge clk);
#1;data_in = testData5[7793];
@(posedge clk);
#1;data_in = testData5[7794];
@(posedge clk);
#1;data_in = testData5[7795];
@(posedge clk);
#1;data_in = testData5[7796];
@(posedge clk);
#1;data_in = testData5[7797];
@(posedge clk);
#1;data_in = testData5[7798];
@(posedge clk);
#1;data_in = testData5[7799];
@(posedge clk);
#1;data_in = testData5[7800];
@(posedge clk);
#1;data_in = testData5[7801];
@(posedge clk);
#1;data_in = testData5[7802];
@(posedge clk);
#1;data_in = testData5[7803];
@(posedge clk);
#1;data_in = testData5[7804];
@(posedge clk);
#1;data_in = testData5[7805];
@(posedge clk);
#1;data_in = testData5[7806];
@(posedge clk);
#1;data_in = testData5[7807];
@(posedge clk);
#1;data_in = testData5[7808];
@(posedge clk);
#1;data_in = testData5[7809];
@(posedge clk);
#1;data_in = testData5[7810];
@(posedge clk);
#1;data_in = testData5[7811];
@(posedge clk);
#1;data_in = testData5[7812];
@(posedge clk);
#1;data_in = testData5[7813];
@(posedge clk);
#1;data_in = testData5[7814];
@(posedge clk);
#1;data_in = testData5[7815];
@(posedge clk);
#1;data_in = testData5[7816];
@(posedge clk);
#1;data_in = testData5[7817];
@(posedge clk);
#1;data_in = testData5[7818];
@(posedge clk);
#1;data_in = testData5[7819];
@(posedge clk);
#1;data_in = testData5[7820];
@(posedge clk);
#1;data_in = testData5[7821];
@(posedge clk);
#1;data_in = testData5[7822];
@(posedge clk);
#1;data_in = testData5[7823];
@(posedge clk);
#1;data_in = testData5[7824];
@(posedge clk);
#1;data_in = testData5[7825];
@(posedge clk);
#1;data_in = testData5[7826];
@(posedge clk);
#1;data_in = testData5[7827];
@(posedge clk);
#1;data_in = testData5[7828];
@(posedge clk);
#1;data_in = testData5[7829];
@(posedge clk);
#1;data_in = testData5[7830];
@(posedge clk);
#1;data_in = testData5[7831];
@(posedge clk);
#1;data_in = testData5[7832];
@(posedge clk);
#1;data_in = testData5[7833];
@(posedge clk);
#1;data_in = testData5[7834];
@(posedge clk);
#1;data_in = testData5[7835];
@(posedge clk);
#1;data_in = testData5[7836];
@(posedge clk);
#1;data_in = testData5[7837];
@(posedge clk);
#1;data_in = testData5[7838];
@(posedge clk);
#1;data_in = testData5[7839];
@(posedge clk);
#1;data_in = testData5[7840];
@(posedge clk);
#1;data_in = testData5[7841];
@(posedge clk);
#1;data_in = testData5[7842];
@(posedge clk);
#1;data_in = testData5[7843];
@(posedge clk);
#1;data_in = testData5[7844];
@(posedge clk);
#1;data_in = testData5[7845];
@(posedge clk);
#1;data_in = testData5[7846];
@(posedge clk);
#1;data_in = testData5[7847];
@(posedge clk);
#1;data_in = testData5[7848];
@(posedge clk);
#1;data_in = testData5[7849];
@(posedge clk);
#1;data_in = testData5[7850];
@(posedge clk);
#1;data_in = testData5[7851];
@(posedge clk);
#1;data_in = testData5[7852];
@(posedge clk);
#1;data_in = testData5[7853];
@(posedge clk);
#1;data_in = testData5[7854];
@(posedge clk);
#1;data_in = testData5[7855];
@(posedge clk);
#1;data_in = testData5[7856];
@(posedge clk);
#1;data_in = testData5[7857];
@(posedge clk);
#1;data_in = testData5[7858];
@(posedge clk);
#1;data_in = testData5[7859];
@(posedge clk);
#1;data_in = testData5[7860];
@(posedge clk);
#1;data_in = testData5[7861];
@(posedge clk);
#1;data_in = testData5[7862];
@(posedge clk);
#1;data_in = testData5[7863];
@(posedge clk);
#1;data_in = testData5[7864];
@(posedge clk);
#1;data_in = testData5[7865];
@(posedge clk);
#1;data_in = testData5[7866];
@(posedge clk);
#1;data_in = testData5[7867];
@(posedge clk);
#1;data_in = testData5[7868];
@(posedge clk);
#1;data_in = testData5[7869];
@(posedge clk);
#1;data_in = testData5[7870];
@(posedge clk);
#1;data_in = testData5[7871];
@(posedge clk);
#1;data_in = testData5[7872];
@(posedge clk);
#1;data_in = testData5[7873];
@(posedge clk);
#1;data_in = testData5[7874];
@(posedge clk);
#1;data_in = testData5[7875];
@(posedge clk);
#1;data_in = testData5[7876];
@(posedge clk);
#1;data_in = testData5[7877];
@(posedge clk);
#1;data_in = testData5[7878];
@(posedge clk);
#1;data_in = testData5[7879];
@(posedge clk);
#1;data_in = testData5[7880];
@(posedge clk);
#1;data_in = testData5[7881];
@(posedge clk);
#1;data_in = testData5[7882];
@(posedge clk);
#1;data_in = testData5[7883];
@(posedge clk);
#1;data_in = testData5[7884];
@(posedge clk);
#1;data_in = testData5[7885];
@(posedge clk);
#1;data_in = testData5[7886];
@(posedge clk);
#1;data_in = testData5[7887];
@(posedge clk);
#1;data_in = testData5[7888];
@(posedge clk);
#1;data_in = testData5[7889];
@(posedge clk);
#1;data_in = testData5[7890];
@(posedge clk);
#1;data_in = testData5[7891];
@(posedge clk);
#1;data_in = testData5[7892];
@(posedge clk);
#1;data_in = testData5[7893];
@(posedge clk);
#1;data_in = testData5[7894];
@(posedge clk);
#1;data_in = testData5[7895];
@(posedge clk);
#1;data_in = testData5[7896];
@(posedge clk);
#1;data_in = testData5[7897];
@(posedge clk);
#1;data_in = testData5[7898];
@(posedge clk);
#1;data_in = testData5[7899];
@(posedge clk);
#1;data_in = testData5[7900];
@(posedge clk);
#1;data_in = testData5[7901];
@(posedge clk);
#1;data_in = testData5[7902];
@(posedge clk);
#1;data_in = testData5[7903];
@(posedge clk);
#1;data_in = testData5[7904];
@(posedge clk);
#1;data_in = testData5[7905];
@(posedge clk);
#1;data_in = testData5[7906];
@(posedge clk);
#1;data_in = testData5[7907];
@(posedge clk);
#1;data_in = testData5[7908];
@(posedge clk);
#1;data_in = testData5[7909];
@(posedge clk);
#1;data_in = testData5[7910];
@(posedge clk);
#1;data_in = testData5[7911];
@(posedge clk);
#1;data_in = testData5[7912];
@(posedge clk);
#1;data_in = testData5[7913];
@(posedge clk);
#1;data_in = testData5[7914];
@(posedge clk);
#1;data_in = testData5[7915];
@(posedge clk);
#1;data_in = testData5[7916];
@(posedge clk);
#1;data_in = testData5[7917];
@(posedge clk);
#1;data_in = testData5[7918];
@(posedge clk);
#1;data_in = testData5[7919];
@(posedge clk);
#1;data_in = testData5[7920];
@(posedge clk);
#1;data_in = testData5[7921];
@(posedge clk);
#1;data_in = testData5[7922];
@(posedge clk);
#1;data_in = testData5[7923];
@(posedge clk);
#1;data_in = testData5[7924];
@(posedge clk);
#1;data_in = testData5[7925];
@(posedge clk);
#1;data_in = testData5[7926];
@(posedge clk);
#1;data_in = testData5[7927];
@(posedge clk);
#1;data_in = testData5[7928];
@(posedge clk);
#1;data_in = testData5[7929];
@(posedge clk);
#1;data_in = testData5[7930];
@(posedge clk);
#1;data_in = testData5[7931];
@(posedge clk);
#1;data_in = testData5[7932];
@(posedge clk);
#1;data_in = testData5[7933];
@(posedge clk);
#1;data_in = testData5[7934];
@(posedge clk);
#1;data_in = testData5[7935];
@(posedge clk);
#1;data_in = testData5[7936];
@(posedge clk);
#1;data_in = testData5[7937];
@(posedge clk);
#1;data_in = testData5[7938];
@(posedge clk);
#1;data_in = testData5[7939];
@(posedge clk);
#1;data_in = testData5[7940];
@(posedge clk);
#1;data_in = testData5[7941];
@(posedge clk);
#1;data_in = testData5[7942];
@(posedge clk);
#1;data_in = testData5[7943];
@(posedge clk);
#1;data_in = testData5[7944];
@(posedge clk);
#1;data_in = testData5[7945];
@(posedge clk);
#1;data_in = testData5[7946];
@(posedge clk);
#1;data_in = testData5[7947];
@(posedge clk);
#1;data_in = testData5[7948];
@(posedge clk);
#1;data_in = testData5[7949];
@(posedge clk);
#1;data_in = testData5[7950];
@(posedge clk);
#1;data_in = testData5[7951];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[7952]; 
@(posedge clk);
#1;data_in = testData5[7953];
@(posedge clk);
#1;data_in = testData5[7954];
@(posedge clk);
#1;data_in = testData5[7955];
@(posedge clk);
#1;data_in = testData5[7956];
@(posedge clk);
#1;data_in = testData5[7957];
@(posedge clk);
#1;data_in = testData5[7958];
@(posedge clk);
#1;data_in = testData5[7959];
@(posedge clk);
#1;data_in = testData5[7960];
@(posedge clk);
#1;data_in = testData5[7961];
@(posedge clk);
#1;data_in = testData5[7962];
@(posedge clk);
#1;data_in = testData5[7963];
@(posedge clk);
#1;data_in = testData5[7964];
@(posedge clk);
#1;data_in = testData5[7965];
@(posedge clk);
#1;data_in = testData5[7966];
@(posedge clk);
#1;data_in = testData5[7967];
@(posedge clk);
#1;data_in = testData5[7968];
@(posedge clk);
#1;data_in = testData5[7969];
@(posedge clk);
#1;data_in = testData5[7970];
@(posedge clk);
#1;data_in = testData5[7971];
@(posedge clk);
#1;data_in = testData5[7972];
@(posedge clk);
#1;data_in = testData5[7973];
@(posedge clk);
#1;data_in = testData5[7974];
@(posedge clk);
#1;data_in = testData5[7975];
@(posedge clk);
#1;data_in = testData5[7976];
@(posedge clk);
#1;data_in = testData5[7977];
@(posedge clk);
#1;data_in = testData5[7978];
@(posedge clk);
#1;data_in = testData5[7979];
@(posedge clk);
#1;data_in = testData5[7980];
@(posedge clk);
#1;data_in = testData5[7981];
@(posedge clk);
#1;data_in = testData5[7982];
@(posedge clk);
#1;data_in = testData5[7983];
@(posedge clk);
#1;data_in = testData5[7984];
@(posedge clk);
#1;data_in = testData5[7985];
@(posedge clk);
#1;data_in = testData5[7986];
@(posedge clk);
#1;data_in = testData5[7987];
@(posedge clk);
#1;data_in = testData5[7988];
@(posedge clk);
#1;data_in = testData5[7989];
@(posedge clk);
#1;data_in = testData5[7990];
@(posedge clk);
#1;data_in = testData5[7991];
@(posedge clk);
#1;data_in = testData5[7992];
@(posedge clk);
#1;data_in = testData5[7993];
@(posedge clk);
#1;data_in = testData5[7994];
@(posedge clk);
#1;data_in = testData5[7995];
@(posedge clk);
#1;data_in = testData5[7996];
@(posedge clk);
#1;data_in = testData5[7997];
@(posedge clk);
#1;data_in = testData5[7998];
@(posedge clk);
#1;data_in = testData5[7999];
@(posedge clk);
#1;data_in = testData5[8000];
@(posedge clk);
#1;data_in = testData5[8001];
@(posedge clk);
#1;data_in = testData5[8002];
@(posedge clk);
#1;data_in = testData5[8003];
@(posedge clk);
#1;data_in = testData5[8004];
@(posedge clk);
#1;data_in = testData5[8005];
@(posedge clk);
#1;data_in = testData5[8006];
@(posedge clk);
#1;data_in = testData5[8007];
@(posedge clk);
#1;data_in = testData5[8008];
@(posedge clk);
#1;data_in = testData5[8009];
@(posedge clk);
#1;data_in = testData5[8010];
@(posedge clk);
#1;data_in = testData5[8011];
@(posedge clk);
#1;data_in = testData5[8012];
@(posedge clk);
#1;data_in = testData5[8013];
@(posedge clk);
#1;data_in = testData5[8014];
@(posedge clk);
#1;data_in = testData5[8015];
@(posedge clk);
#1;data_in = testData5[8016];
@(posedge clk);
#1;data_in = testData5[8017];
@(posedge clk);
#1;data_in = testData5[8018];
@(posedge clk);
#1;data_in = testData5[8019];
@(posedge clk);
#1;data_in = testData5[8020];
@(posedge clk);
#1;data_in = testData5[8021];
@(posedge clk);
#1;data_in = testData5[8022];
@(posedge clk);
#1;data_in = testData5[8023];
@(posedge clk);
#1;data_in = testData5[8024];
@(posedge clk);
#1;data_in = testData5[8025];
@(posedge clk);
#1;data_in = testData5[8026];
@(posedge clk);
#1;data_in = testData5[8027];
@(posedge clk);
#1;data_in = testData5[8028];
@(posedge clk);
#1;data_in = testData5[8029];
@(posedge clk);
#1;data_in = testData5[8030];
@(posedge clk);
#1;data_in = testData5[8031];
@(posedge clk);
#1;data_in = testData5[8032];
@(posedge clk);
#1;data_in = testData5[8033];
@(posedge clk);
#1;data_in = testData5[8034];
@(posedge clk);
#1;data_in = testData5[8035];
@(posedge clk);
#1;data_in = testData5[8036];
@(posedge clk);
#1;data_in = testData5[8037];
@(posedge clk);
#1;data_in = testData5[8038];
@(posedge clk);
#1;data_in = testData5[8039];
@(posedge clk);
#1;data_in = testData5[8040];
@(posedge clk);
#1;data_in = testData5[8041];
@(posedge clk);
#1;data_in = testData5[8042];
@(posedge clk);
#1;data_in = testData5[8043];
@(posedge clk);
#1;data_in = testData5[8044];
@(posedge clk);
#1;data_in = testData5[8045];
@(posedge clk);
#1;data_in = testData5[8046];
@(posedge clk);
#1;data_in = testData5[8047];
@(posedge clk);
#1;data_in = testData5[8048];
@(posedge clk);
#1;data_in = testData5[8049];
@(posedge clk);
#1;data_in = testData5[8050];
@(posedge clk);
#1;data_in = testData5[8051];
@(posedge clk);
#1;data_in = testData5[8052];
@(posedge clk);
#1;data_in = testData5[8053];
@(posedge clk);
#1;data_in = testData5[8054];
@(posedge clk);
#1;data_in = testData5[8055];
@(posedge clk);
#1;data_in = testData5[8056];
@(posedge clk);
#1;data_in = testData5[8057];
@(posedge clk);
#1;data_in = testData5[8058];
@(posedge clk);
#1;data_in = testData5[8059];
@(posedge clk);
#1;data_in = testData5[8060];
@(posedge clk);
#1;data_in = testData5[8061];
@(posedge clk);
#1;data_in = testData5[8062];
@(posedge clk);
#1;data_in = testData5[8063];
@(posedge clk);
#1;data_in = testData5[8064];
@(posedge clk);
#1;data_in = testData5[8065];
@(posedge clk);
#1;data_in = testData5[8066];
@(posedge clk);
#1;data_in = testData5[8067];
@(posedge clk);
#1;data_in = testData5[8068];
@(posedge clk);
#1;data_in = testData5[8069];
@(posedge clk);
#1;data_in = testData5[8070];
@(posedge clk);
#1;data_in = testData5[8071];
@(posedge clk);
#1;data_in = testData5[8072];
@(posedge clk);
#1;data_in = testData5[8073];
@(posedge clk);
#1;data_in = testData5[8074];
@(posedge clk);
#1;data_in = testData5[8075];
@(posedge clk);
#1;data_in = testData5[8076];
@(posedge clk);
#1;data_in = testData5[8077];
@(posedge clk);
#1;data_in = testData5[8078];
@(posedge clk);
#1;data_in = testData5[8079];
@(posedge clk);
#1;data_in = testData5[8080];
@(posedge clk);
#1;data_in = testData5[8081];
@(posedge clk);
#1;data_in = testData5[8082];
@(posedge clk);
#1;data_in = testData5[8083];
@(posedge clk);
#1;data_in = testData5[8084];
@(posedge clk);
#1;data_in = testData5[8085];
@(posedge clk);
#1;data_in = testData5[8086];
@(posedge clk);
#1;data_in = testData5[8087];
@(posedge clk);
#1;data_in = testData5[8088];
@(posedge clk);
#1;data_in = testData5[8089];
@(posedge clk);
#1;data_in = testData5[8090];
@(posedge clk);
#1;data_in = testData5[8091];
@(posedge clk);
#1;data_in = testData5[8092];
@(posedge clk);
#1;data_in = testData5[8093];
@(posedge clk);
#1;data_in = testData5[8094];
@(posedge clk);
#1;data_in = testData5[8095];
@(posedge clk);
#1;data_in = testData5[8096];
@(posedge clk);
#1;data_in = testData5[8097];
@(posedge clk);
#1;data_in = testData5[8098];
@(posedge clk);
#1;data_in = testData5[8099];
@(posedge clk);
#1;data_in = testData5[8100];
@(posedge clk);
#1;data_in = testData5[8101];
@(posedge clk);
#1;data_in = testData5[8102];
@(posedge clk);
#1;data_in = testData5[8103];
@(posedge clk);
#1;data_in = testData5[8104];
@(posedge clk);
#1;data_in = testData5[8105];
@(posedge clk);
#1;data_in = testData5[8106];
@(posedge clk);
#1;data_in = testData5[8107];
@(posedge clk);
#1;data_in = testData5[8108];
@(posedge clk);
#1;data_in = testData5[8109];
@(posedge clk);
#1;data_in = testData5[8110];
@(posedge clk);
#1;data_in = testData5[8111];
@(posedge clk);
#1;data_in = testData5[8112];
@(posedge clk);
#1;data_in = testData5[8113];
@(posedge clk);
#1;data_in = testData5[8114];
@(posedge clk);
#1;data_in = testData5[8115];
@(posedge clk);
#1;data_in = testData5[8116];
@(posedge clk);
#1;data_in = testData5[8117];
@(posedge clk);
#1;data_in = testData5[8118];
@(posedge clk);
#1;data_in = testData5[8119];
@(posedge clk);
#1;data_in = testData5[8120];
@(posedge clk);
#1;data_in = testData5[8121];
@(posedge clk);
#1;data_in = testData5[8122];
@(posedge clk);
#1;data_in = testData5[8123];
@(posedge clk);
#1;data_in = testData5[8124];
@(posedge clk);
#1;data_in = testData5[8125];
@(posedge clk);
#1;data_in = testData5[8126];
@(posedge clk);
#1;data_in = testData5[8127];
@(posedge clk);
#1;data_in = testData5[8128];
@(posedge clk);
#1;data_in = testData5[8129];
@(posedge clk);
#1;data_in = testData5[8130];
@(posedge clk);
#1;data_in = testData5[8131];
@(posedge clk);
#1;data_in = testData5[8132];
@(posedge clk);
#1;data_in = testData5[8133];
@(posedge clk);
#1;data_in = testData5[8134];
@(posedge clk);
#1;data_in = testData5[8135];
@(posedge clk);
#1;data_in = testData5[8136];
@(posedge clk);
#1;data_in = testData5[8137];
@(posedge clk);
#1;data_in = testData5[8138];
@(posedge clk);
#1;data_in = testData5[8139];
@(posedge clk);
#1;data_in = testData5[8140];
@(posedge clk);
#1;data_in = testData5[8141];
@(posedge clk);
#1;data_in = testData5[8142];
@(posedge clk);
#1;data_in = testData5[8143];
@(posedge clk);
#1;data_in = testData5[8144];
@(posedge clk);
#1;data_in = testData5[8145];
@(posedge clk);
#1;data_in = testData5[8146];
@(posedge clk);
#1;data_in = testData5[8147];
@(posedge clk);
#1;data_in = testData5[8148];
@(posedge clk);
#1;data_in = testData5[8149];
@(posedge clk);
#1;data_in = testData5[8150];
@(posedge clk);
#1;data_in = testData5[8151];
@(posedge clk);
#1;data_in = testData5[8152];
@(posedge clk);
#1;data_in = testData5[8153];
@(posedge clk);
#1;data_in = testData5[8154];
@(posedge clk);
#1;data_in = testData5[8155];
@(posedge clk);
#1;data_in = testData5[8156];
@(posedge clk);
#1;data_in = testData5[8157];
@(posedge clk);
#1;data_in = testData5[8158];
@(posedge clk);
#1;data_in = testData5[8159];
@(posedge clk);
#1;data_in = testData5[8160];
@(posedge clk);
#1;data_in = testData5[8161];
@(posedge clk);
#1;data_in = testData5[8162];
@(posedge clk);
#1;data_in = testData5[8163];
@(posedge clk);
#1;data_in = testData5[8164];
@(posedge clk);
#1;data_in = testData5[8165];
@(posedge clk);
#1;data_in = testData5[8166];
@(posedge clk);
#1;data_in = testData5[8167];
@(posedge clk);
#1;data_in = testData5[8168];
@(posedge clk);
#1;data_in = testData5[8169];
@(posedge clk);
#1;data_in = testData5[8170];
@(posedge clk);
#1;data_in = testData5[8171];
@(posedge clk);
#1;data_in = testData5[8172];
@(posedge clk);
#1;data_in = testData5[8173];
@(posedge clk);
#1;data_in = testData5[8174];
@(posedge clk);
#1;data_in = testData5[8175];
@(posedge clk);
#1;data_in = testData5[8176];
@(posedge clk);
#1;data_in = testData5[8177];
@(posedge clk);
#1;data_in = testData5[8178];
@(posedge clk);
#1;data_in = testData5[8179];
@(posedge clk);
#1;data_in = testData5[8180];
@(posedge clk);
#1;data_in = testData5[8181];
@(posedge clk);
#1;data_in = testData5[8182];
@(posedge clk);
#1;data_in = testData5[8183];
@(posedge clk);
#1;data_in = testData5[8184];
@(posedge clk);
#1;data_in = testData5[8185];
@(posedge clk);
#1;data_in = testData5[8186];
@(posedge clk);
#1;data_in = testData5[8187];
@(posedge clk);
#1;data_in = testData5[8188];
@(posedge clk);
#1;data_in = testData5[8189];
@(posedge clk);
#1;data_in = testData5[8190];
@(posedge clk);
#1;data_in = testData5[8191];
@(posedge clk);
#1;data_in = testData5[8192];
@(posedge clk);
#1;data_in = testData5[8193];
@(posedge clk);
#1;data_in = testData5[8194];
@(posedge clk);
#1;data_in = testData5[8195];
@(posedge clk);
#1;data_in = testData5[8196];
@(posedge clk);
#1;data_in = testData5[8197];
@(posedge clk);
#1;data_in = testData5[8198];
@(posedge clk);
#1;data_in = testData5[8199];
@(posedge clk);
#1;data_in = testData5[8200];
@(posedge clk);
#1;data_in = testData5[8201];
@(posedge clk);
#1;data_in = testData5[8202];
@(posedge clk);
#1;data_in = testData5[8203];
@(posedge clk);
#1;data_in = testData5[8204];
@(posedge clk);
#1;data_in = testData5[8205];
@(posedge clk);
#1;data_in = testData5[8206];
@(posedge clk);
#1;data_in = testData5[8207];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[8208]; 
@(posedge clk);
#1;data_in = testData5[8209];
@(posedge clk);
#1;data_in = testData5[8210];
@(posedge clk);
#1;data_in = testData5[8211];
@(posedge clk);
#1;data_in = testData5[8212];
@(posedge clk);
#1;data_in = testData5[8213];
@(posedge clk);
#1;data_in = testData5[8214];
@(posedge clk);
#1;data_in = testData5[8215];
@(posedge clk);
#1;data_in = testData5[8216];
@(posedge clk);
#1;data_in = testData5[8217];
@(posedge clk);
#1;data_in = testData5[8218];
@(posedge clk);
#1;data_in = testData5[8219];
@(posedge clk);
#1;data_in = testData5[8220];
@(posedge clk);
#1;data_in = testData5[8221];
@(posedge clk);
#1;data_in = testData5[8222];
@(posedge clk);
#1;data_in = testData5[8223];
@(posedge clk);
#1;data_in = testData5[8224];
@(posedge clk);
#1;data_in = testData5[8225];
@(posedge clk);
#1;data_in = testData5[8226];
@(posedge clk);
#1;data_in = testData5[8227];
@(posedge clk);
#1;data_in = testData5[8228];
@(posedge clk);
#1;data_in = testData5[8229];
@(posedge clk);
#1;data_in = testData5[8230];
@(posedge clk);
#1;data_in = testData5[8231];
@(posedge clk);
#1;data_in = testData5[8232];
@(posedge clk);
#1;data_in = testData5[8233];
@(posedge clk);
#1;data_in = testData5[8234];
@(posedge clk);
#1;data_in = testData5[8235];
@(posedge clk);
#1;data_in = testData5[8236];
@(posedge clk);
#1;data_in = testData5[8237];
@(posedge clk);
#1;data_in = testData5[8238];
@(posedge clk);
#1;data_in = testData5[8239];
@(posedge clk);
#1;data_in = testData5[8240];
@(posedge clk);
#1;data_in = testData5[8241];
@(posedge clk);
#1;data_in = testData5[8242];
@(posedge clk);
#1;data_in = testData5[8243];
@(posedge clk);
#1;data_in = testData5[8244];
@(posedge clk);
#1;data_in = testData5[8245];
@(posedge clk);
#1;data_in = testData5[8246];
@(posedge clk);
#1;data_in = testData5[8247];
@(posedge clk);
#1;data_in = testData5[8248];
@(posedge clk);
#1;data_in = testData5[8249];
@(posedge clk);
#1;data_in = testData5[8250];
@(posedge clk);
#1;data_in = testData5[8251];
@(posedge clk);
#1;data_in = testData5[8252];
@(posedge clk);
#1;data_in = testData5[8253];
@(posedge clk);
#1;data_in = testData5[8254];
@(posedge clk);
#1;data_in = testData5[8255];
@(posedge clk);
#1;data_in = testData5[8256];
@(posedge clk);
#1;data_in = testData5[8257];
@(posedge clk);
#1;data_in = testData5[8258];
@(posedge clk);
#1;data_in = testData5[8259];
@(posedge clk);
#1;data_in = testData5[8260];
@(posedge clk);
#1;data_in = testData5[8261];
@(posedge clk);
#1;data_in = testData5[8262];
@(posedge clk);
#1;data_in = testData5[8263];
@(posedge clk);
#1;data_in = testData5[8264];
@(posedge clk);
#1;data_in = testData5[8265];
@(posedge clk);
#1;data_in = testData5[8266];
@(posedge clk);
#1;data_in = testData5[8267];
@(posedge clk);
#1;data_in = testData5[8268];
@(posedge clk);
#1;data_in = testData5[8269];
@(posedge clk);
#1;data_in = testData5[8270];
@(posedge clk);
#1;data_in = testData5[8271];
@(posedge clk);
#1;data_in = testData5[8272];
@(posedge clk);
#1;data_in = testData5[8273];
@(posedge clk);
#1;data_in = testData5[8274];
@(posedge clk);
#1;data_in = testData5[8275];
@(posedge clk);
#1;data_in = testData5[8276];
@(posedge clk);
#1;data_in = testData5[8277];
@(posedge clk);
#1;data_in = testData5[8278];
@(posedge clk);
#1;data_in = testData5[8279];
@(posedge clk);
#1;data_in = testData5[8280];
@(posedge clk);
#1;data_in = testData5[8281];
@(posedge clk);
#1;data_in = testData5[8282];
@(posedge clk);
#1;data_in = testData5[8283];
@(posedge clk);
#1;data_in = testData5[8284];
@(posedge clk);
#1;data_in = testData5[8285];
@(posedge clk);
#1;data_in = testData5[8286];
@(posedge clk);
#1;data_in = testData5[8287];
@(posedge clk);
#1;data_in = testData5[8288];
@(posedge clk);
#1;data_in = testData5[8289];
@(posedge clk);
#1;data_in = testData5[8290];
@(posedge clk);
#1;data_in = testData5[8291];
@(posedge clk);
#1;data_in = testData5[8292];
@(posedge clk);
#1;data_in = testData5[8293];
@(posedge clk);
#1;data_in = testData5[8294];
@(posedge clk);
#1;data_in = testData5[8295];
@(posedge clk);
#1;data_in = testData5[8296];
@(posedge clk);
#1;data_in = testData5[8297];
@(posedge clk);
#1;data_in = testData5[8298];
@(posedge clk);
#1;data_in = testData5[8299];
@(posedge clk);
#1;data_in = testData5[8300];
@(posedge clk);
#1;data_in = testData5[8301];
@(posedge clk);
#1;data_in = testData5[8302];
@(posedge clk);
#1;data_in = testData5[8303];
@(posedge clk);
#1;data_in = testData5[8304];
@(posedge clk);
#1;data_in = testData5[8305];
@(posedge clk);
#1;data_in = testData5[8306];
@(posedge clk);
#1;data_in = testData5[8307];
@(posedge clk);
#1;data_in = testData5[8308];
@(posedge clk);
#1;data_in = testData5[8309];
@(posedge clk);
#1;data_in = testData5[8310];
@(posedge clk);
#1;data_in = testData5[8311];
@(posedge clk);
#1;data_in = testData5[8312];
@(posedge clk);
#1;data_in = testData5[8313];
@(posedge clk);
#1;data_in = testData5[8314];
@(posedge clk);
#1;data_in = testData5[8315];
@(posedge clk);
#1;data_in = testData5[8316];
@(posedge clk);
#1;data_in = testData5[8317];
@(posedge clk);
#1;data_in = testData5[8318];
@(posedge clk);
#1;data_in = testData5[8319];
@(posedge clk);
#1;data_in = testData5[8320];
@(posedge clk);
#1;data_in = testData5[8321];
@(posedge clk);
#1;data_in = testData5[8322];
@(posedge clk);
#1;data_in = testData5[8323];
@(posedge clk);
#1;data_in = testData5[8324];
@(posedge clk);
#1;data_in = testData5[8325];
@(posedge clk);
#1;data_in = testData5[8326];
@(posedge clk);
#1;data_in = testData5[8327];
@(posedge clk);
#1;data_in = testData5[8328];
@(posedge clk);
#1;data_in = testData5[8329];
@(posedge clk);
#1;data_in = testData5[8330];
@(posedge clk);
#1;data_in = testData5[8331];
@(posedge clk);
#1;data_in = testData5[8332];
@(posedge clk);
#1;data_in = testData5[8333];
@(posedge clk);
#1;data_in = testData5[8334];
@(posedge clk);
#1;data_in = testData5[8335];
@(posedge clk);
#1;data_in = testData5[8336];
@(posedge clk);
#1;data_in = testData5[8337];
@(posedge clk);
#1;data_in = testData5[8338];
@(posedge clk);
#1;data_in = testData5[8339];
@(posedge clk);
#1;data_in = testData5[8340];
@(posedge clk);
#1;data_in = testData5[8341];
@(posedge clk);
#1;data_in = testData5[8342];
@(posedge clk);
#1;data_in = testData5[8343];
@(posedge clk);
#1;data_in = testData5[8344];
@(posedge clk);
#1;data_in = testData5[8345];
@(posedge clk);
#1;data_in = testData5[8346];
@(posedge clk);
#1;data_in = testData5[8347];
@(posedge clk);
#1;data_in = testData5[8348];
@(posedge clk);
#1;data_in = testData5[8349];
@(posedge clk);
#1;data_in = testData5[8350];
@(posedge clk);
#1;data_in = testData5[8351];
@(posedge clk);
#1;data_in = testData5[8352];
@(posedge clk);
#1;data_in = testData5[8353];
@(posedge clk);
#1;data_in = testData5[8354];
@(posedge clk);
#1;data_in = testData5[8355];
@(posedge clk);
#1;data_in = testData5[8356];
@(posedge clk);
#1;data_in = testData5[8357];
@(posedge clk);
#1;data_in = testData5[8358];
@(posedge clk);
#1;data_in = testData5[8359];
@(posedge clk);
#1;data_in = testData5[8360];
@(posedge clk);
#1;data_in = testData5[8361];
@(posedge clk);
#1;data_in = testData5[8362];
@(posedge clk);
#1;data_in = testData5[8363];
@(posedge clk);
#1;data_in = testData5[8364];
@(posedge clk);
#1;data_in = testData5[8365];
@(posedge clk);
#1;data_in = testData5[8366];
@(posedge clk);
#1;data_in = testData5[8367];
@(posedge clk);
#1;data_in = testData5[8368];
@(posedge clk);
#1;data_in = testData5[8369];
@(posedge clk);
#1;data_in = testData5[8370];
@(posedge clk);
#1;data_in = testData5[8371];
@(posedge clk);
#1;data_in = testData5[8372];
@(posedge clk);
#1;data_in = testData5[8373];
@(posedge clk);
#1;data_in = testData5[8374];
@(posedge clk);
#1;data_in = testData5[8375];
@(posedge clk);
#1;data_in = testData5[8376];
@(posedge clk);
#1;data_in = testData5[8377];
@(posedge clk);
#1;data_in = testData5[8378];
@(posedge clk);
#1;data_in = testData5[8379];
@(posedge clk);
#1;data_in = testData5[8380];
@(posedge clk);
#1;data_in = testData5[8381];
@(posedge clk);
#1;data_in = testData5[8382];
@(posedge clk);
#1;data_in = testData5[8383];
@(posedge clk);
#1;data_in = testData5[8384];
@(posedge clk);
#1;data_in = testData5[8385];
@(posedge clk);
#1;data_in = testData5[8386];
@(posedge clk);
#1;data_in = testData5[8387];
@(posedge clk);
#1;data_in = testData5[8388];
@(posedge clk);
#1;data_in = testData5[8389];
@(posedge clk);
#1;data_in = testData5[8390];
@(posedge clk);
#1;data_in = testData5[8391];
@(posedge clk);
#1;data_in = testData5[8392];
@(posedge clk);
#1;data_in = testData5[8393];
@(posedge clk);
#1;data_in = testData5[8394];
@(posedge clk);
#1;data_in = testData5[8395];
@(posedge clk);
#1;data_in = testData5[8396];
@(posedge clk);
#1;data_in = testData5[8397];
@(posedge clk);
#1;data_in = testData5[8398];
@(posedge clk);
#1;data_in = testData5[8399];
@(posedge clk);
#1;data_in = testData5[8400];
@(posedge clk);
#1;data_in = testData5[8401];
@(posedge clk);
#1;data_in = testData5[8402];
@(posedge clk);
#1;data_in = testData5[8403];
@(posedge clk);
#1;data_in = testData5[8404];
@(posedge clk);
#1;data_in = testData5[8405];
@(posedge clk);
#1;data_in = testData5[8406];
@(posedge clk);
#1;data_in = testData5[8407];
@(posedge clk);
#1;data_in = testData5[8408];
@(posedge clk);
#1;data_in = testData5[8409];
@(posedge clk);
#1;data_in = testData5[8410];
@(posedge clk);
#1;data_in = testData5[8411];
@(posedge clk);
#1;data_in = testData5[8412];
@(posedge clk);
#1;data_in = testData5[8413];
@(posedge clk);
#1;data_in = testData5[8414];
@(posedge clk);
#1;data_in = testData5[8415];
@(posedge clk);
#1;data_in = testData5[8416];
@(posedge clk);
#1;data_in = testData5[8417];
@(posedge clk);
#1;data_in = testData5[8418];
@(posedge clk);
#1;data_in = testData5[8419];
@(posedge clk);
#1;data_in = testData5[8420];
@(posedge clk);
#1;data_in = testData5[8421];
@(posedge clk);
#1;data_in = testData5[8422];
@(posedge clk);
#1;data_in = testData5[8423];
@(posedge clk);
#1;data_in = testData5[8424];
@(posedge clk);
#1;data_in = testData5[8425];
@(posedge clk);
#1;data_in = testData5[8426];
@(posedge clk);
#1;data_in = testData5[8427];
@(posedge clk);
#1;data_in = testData5[8428];
@(posedge clk);
#1;data_in = testData5[8429];
@(posedge clk);
#1;data_in = testData5[8430];
@(posedge clk);
#1;data_in = testData5[8431];
@(posedge clk);
#1;data_in = testData5[8432];
@(posedge clk);
#1;data_in = testData5[8433];
@(posedge clk);
#1;data_in = testData5[8434];
@(posedge clk);
#1;data_in = testData5[8435];
@(posedge clk);
#1;data_in = testData5[8436];
@(posedge clk);
#1;data_in = testData5[8437];
@(posedge clk);
#1;data_in = testData5[8438];
@(posedge clk);
#1;data_in = testData5[8439];
@(posedge clk);
#1;data_in = testData5[8440];
@(posedge clk);
#1;data_in = testData5[8441];
@(posedge clk);
#1;data_in = testData5[8442];
@(posedge clk);
#1;data_in = testData5[8443];
@(posedge clk);
#1;data_in = testData5[8444];
@(posedge clk);
#1;data_in = testData5[8445];
@(posedge clk);
#1;data_in = testData5[8446];
@(posedge clk);
#1;data_in = testData5[8447];
@(posedge clk);
#1;data_in = testData5[8448];
@(posedge clk);
#1;data_in = testData5[8449];
@(posedge clk);
#1;data_in = testData5[8450];
@(posedge clk);
#1;data_in = testData5[8451];
@(posedge clk);
#1;data_in = testData5[8452];
@(posedge clk);
#1;data_in = testData5[8453];
@(posedge clk);
#1;data_in = testData5[8454];
@(posedge clk);
#1;data_in = testData5[8455];
@(posedge clk);
#1;data_in = testData5[8456];
@(posedge clk);
#1;data_in = testData5[8457];
@(posedge clk);
#1;data_in = testData5[8458];
@(posedge clk);
#1;data_in = testData5[8459];
@(posedge clk);
#1;data_in = testData5[8460];
@(posedge clk);
#1;data_in = testData5[8461];
@(posedge clk);
#1;data_in = testData5[8462];
@(posedge clk);
#1;data_in = testData5[8463];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[8464]; 
@(posedge clk);
#1;data_in = testData5[8465];
@(posedge clk);
#1;data_in = testData5[8466];
@(posedge clk);
#1;data_in = testData5[8467];
@(posedge clk);
#1;data_in = testData5[8468];
@(posedge clk);
#1;data_in = testData5[8469];
@(posedge clk);
#1;data_in = testData5[8470];
@(posedge clk);
#1;data_in = testData5[8471];
@(posedge clk);
#1;data_in = testData5[8472];
@(posedge clk);
#1;data_in = testData5[8473];
@(posedge clk);
#1;data_in = testData5[8474];
@(posedge clk);
#1;data_in = testData5[8475];
@(posedge clk);
#1;data_in = testData5[8476];
@(posedge clk);
#1;data_in = testData5[8477];
@(posedge clk);
#1;data_in = testData5[8478];
@(posedge clk);
#1;data_in = testData5[8479];
@(posedge clk);
#1;data_in = testData5[8480];
@(posedge clk);
#1;data_in = testData5[8481];
@(posedge clk);
#1;data_in = testData5[8482];
@(posedge clk);
#1;data_in = testData5[8483];
@(posedge clk);
#1;data_in = testData5[8484];
@(posedge clk);
#1;data_in = testData5[8485];
@(posedge clk);
#1;data_in = testData5[8486];
@(posedge clk);
#1;data_in = testData5[8487];
@(posedge clk);
#1;data_in = testData5[8488];
@(posedge clk);
#1;data_in = testData5[8489];
@(posedge clk);
#1;data_in = testData5[8490];
@(posedge clk);
#1;data_in = testData5[8491];
@(posedge clk);
#1;data_in = testData5[8492];
@(posedge clk);
#1;data_in = testData5[8493];
@(posedge clk);
#1;data_in = testData5[8494];
@(posedge clk);
#1;data_in = testData5[8495];
@(posedge clk);
#1;data_in = testData5[8496];
@(posedge clk);
#1;data_in = testData5[8497];
@(posedge clk);
#1;data_in = testData5[8498];
@(posedge clk);
#1;data_in = testData5[8499];
@(posedge clk);
#1;data_in = testData5[8500];
@(posedge clk);
#1;data_in = testData5[8501];
@(posedge clk);
#1;data_in = testData5[8502];
@(posedge clk);
#1;data_in = testData5[8503];
@(posedge clk);
#1;data_in = testData5[8504];
@(posedge clk);
#1;data_in = testData5[8505];
@(posedge clk);
#1;data_in = testData5[8506];
@(posedge clk);
#1;data_in = testData5[8507];
@(posedge clk);
#1;data_in = testData5[8508];
@(posedge clk);
#1;data_in = testData5[8509];
@(posedge clk);
#1;data_in = testData5[8510];
@(posedge clk);
#1;data_in = testData5[8511];
@(posedge clk);
#1;data_in = testData5[8512];
@(posedge clk);
#1;data_in = testData5[8513];
@(posedge clk);
#1;data_in = testData5[8514];
@(posedge clk);
#1;data_in = testData5[8515];
@(posedge clk);
#1;data_in = testData5[8516];
@(posedge clk);
#1;data_in = testData5[8517];
@(posedge clk);
#1;data_in = testData5[8518];
@(posedge clk);
#1;data_in = testData5[8519];
@(posedge clk);
#1;data_in = testData5[8520];
@(posedge clk);
#1;data_in = testData5[8521];
@(posedge clk);
#1;data_in = testData5[8522];
@(posedge clk);
#1;data_in = testData5[8523];
@(posedge clk);
#1;data_in = testData5[8524];
@(posedge clk);
#1;data_in = testData5[8525];
@(posedge clk);
#1;data_in = testData5[8526];
@(posedge clk);
#1;data_in = testData5[8527];
@(posedge clk);
#1;data_in = testData5[8528];
@(posedge clk);
#1;data_in = testData5[8529];
@(posedge clk);
#1;data_in = testData5[8530];
@(posedge clk);
#1;data_in = testData5[8531];
@(posedge clk);
#1;data_in = testData5[8532];
@(posedge clk);
#1;data_in = testData5[8533];
@(posedge clk);
#1;data_in = testData5[8534];
@(posedge clk);
#1;data_in = testData5[8535];
@(posedge clk);
#1;data_in = testData5[8536];
@(posedge clk);
#1;data_in = testData5[8537];
@(posedge clk);
#1;data_in = testData5[8538];
@(posedge clk);
#1;data_in = testData5[8539];
@(posedge clk);
#1;data_in = testData5[8540];
@(posedge clk);
#1;data_in = testData5[8541];
@(posedge clk);
#1;data_in = testData5[8542];
@(posedge clk);
#1;data_in = testData5[8543];
@(posedge clk);
#1;data_in = testData5[8544];
@(posedge clk);
#1;data_in = testData5[8545];
@(posedge clk);
#1;data_in = testData5[8546];
@(posedge clk);
#1;data_in = testData5[8547];
@(posedge clk);
#1;data_in = testData5[8548];
@(posedge clk);
#1;data_in = testData5[8549];
@(posedge clk);
#1;data_in = testData5[8550];
@(posedge clk);
#1;data_in = testData5[8551];
@(posedge clk);
#1;data_in = testData5[8552];
@(posedge clk);
#1;data_in = testData5[8553];
@(posedge clk);
#1;data_in = testData5[8554];
@(posedge clk);
#1;data_in = testData5[8555];
@(posedge clk);
#1;data_in = testData5[8556];
@(posedge clk);
#1;data_in = testData5[8557];
@(posedge clk);
#1;data_in = testData5[8558];
@(posedge clk);
#1;data_in = testData5[8559];
@(posedge clk);
#1;data_in = testData5[8560];
@(posedge clk);
#1;data_in = testData5[8561];
@(posedge clk);
#1;data_in = testData5[8562];
@(posedge clk);
#1;data_in = testData5[8563];
@(posedge clk);
#1;data_in = testData5[8564];
@(posedge clk);
#1;data_in = testData5[8565];
@(posedge clk);
#1;data_in = testData5[8566];
@(posedge clk);
#1;data_in = testData5[8567];
@(posedge clk);
#1;data_in = testData5[8568];
@(posedge clk);
#1;data_in = testData5[8569];
@(posedge clk);
#1;data_in = testData5[8570];
@(posedge clk);
#1;data_in = testData5[8571];
@(posedge clk);
#1;data_in = testData5[8572];
@(posedge clk);
#1;data_in = testData5[8573];
@(posedge clk);
#1;data_in = testData5[8574];
@(posedge clk);
#1;data_in = testData5[8575];
@(posedge clk);
#1;data_in = testData5[8576];
@(posedge clk);
#1;data_in = testData5[8577];
@(posedge clk);
#1;data_in = testData5[8578];
@(posedge clk);
#1;data_in = testData5[8579];
@(posedge clk);
#1;data_in = testData5[8580];
@(posedge clk);
#1;data_in = testData5[8581];
@(posedge clk);
#1;data_in = testData5[8582];
@(posedge clk);
#1;data_in = testData5[8583];
@(posedge clk);
#1;data_in = testData5[8584];
@(posedge clk);
#1;data_in = testData5[8585];
@(posedge clk);
#1;data_in = testData5[8586];
@(posedge clk);
#1;data_in = testData5[8587];
@(posedge clk);
#1;data_in = testData5[8588];
@(posedge clk);
#1;data_in = testData5[8589];
@(posedge clk);
#1;data_in = testData5[8590];
@(posedge clk);
#1;data_in = testData5[8591];
@(posedge clk);
#1;data_in = testData5[8592];
@(posedge clk);
#1;data_in = testData5[8593];
@(posedge clk);
#1;data_in = testData5[8594];
@(posedge clk);
#1;data_in = testData5[8595];
@(posedge clk);
#1;data_in = testData5[8596];
@(posedge clk);
#1;data_in = testData5[8597];
@(posedge clk);
#1;data_in = testData5[8598];
@(posedge clk);
#1;data_in = testData5[8599];
@(posedge clk);
#1;data_in = testData5[8600];
@(posedge clk);
#1;data_in = testData5[8601];
@(posedge clk);
#1;data_in = testData5[8602];
@(posedge clk);
#1;data_in = testData5[8603];
@(posedge clk);
#1;data_in = testData5[8604];
@(posedge clk);
#1;data_in = testData5[8605];
@(posedge clk);
#1;data_in = testData5[8606];
@(posedge clk);
#1;data_in = testData5[8607];
@(posedge clk);
#1;data_in = testData5[8608];
@(posedge clk);
#1;data_in = testData5[8609];
@(posedge clk);
#1;data_in = testData5[8610];
@(posedge clk);
#1;data_in = testData5[8611];
@(posedge clk);
#1;data_in = testData5[8612];
@(posedge clk);
#1;data_in = testData5[8613];
@(posedge clk);
#1;data_in = testData5[8614];
@(posedge clk);
#1;data_in = testData5[8615];
@(posedge clk);
#1;data_in = testData5[8616];
@(posedge clk);
#1;data_in = testData5[8617];
@(posedge clk);
#1;data_in = testData5[8618];
@(posedge clk);
#1;data_in = testData5[8619];
@(posedge clk);
#1;data_in = testData5[8620];
@(posedge clk);
#1;data_in = testData5[8621];
@(posedge clk);
#1;data_in = testData5[8622];
@(posedge clk);
#1;data_in = testData5[8623];
@(posedge clk);
#1;data_in = testData5[8624];
@(posedge clk);
#1;data_in = testData5[8625];
@(posedge clk);
#1;data_in = testData5[8626];
@(posedge clk);
#1;data_in = testData5[8627];
@(posedge clk);
#1;data_in = testData5[8628];
@(posedge clk);
#1;data_in = testData5[8629];
@(posedge clk);
#1;data_in = testData5[8630];
@(posedge clk);
#1;data_in = testData5[8631];
@(posedge clk);
#1;data_in = testData5[8632];
@(posedge clk);
#1;data_in = testData5[8633];
@(posedge clk);
#1;data_in = testData5[8634];
@(posedge clk);
#1;data_in = testData5[8635];
@(posedge clk);
#1;data_in = testData5[8636];
@(posedge clk);
#1;data_in = testData5[8637];
@(posedge clk);
#1;data_in = testData5[8638];
@(posedge clk);
#1;data_in = testData5[8639];
@(posedge clk);
#1;data_in = testData5[8640];
@(posedge clk);
#1;data_in = testData5[8641];
@(posedge clk);
#1;data_in = testData5[8642];
@(posedge clk);
#1;data_in = testData5[8643];
@(posedge clk);
#1;data_in = testData5[8644];
@(posedge clk);
#1;data_in = testData5[8645];
@(posedge clk);
#1;data_in = testData5[8646];
@(posedge clk);
#1;data_in = testData5[8647];
@(posedge clk);
#1;data_in = testData5[8648];
@(posedge clk);
#1;data_in = testData5[8649];
@(posedge clk);
#1;data_in = testData5[8650];
@(posedge clk);
#1;data_in = testData5[8651];
@(posedge clk);
#1;data_in = testData5[8652];
@(posedge clk);
#1;data_in = testData5[8653];
@(posedge clk);
#1;data_in = testData5[8654];
@(posedge clk);
#1;data_in = testData5[8655];
@(posedge clk);
#1;data_in = testData5[8656];
@(posedge clk);
#1;data_in = testData5[8657];
@(posedge clk);
#1;data_in = testData5[8658];
@(posedge clk);
#1;data_in = testData5[8659];
@(posedge clk);
#1;data_in = testData5[8660];
@(posedge clk);
#1;data_in = testData5[8661];
@(posedge clk);
#1;data_in = testData5[8662];
@(posedge clk);
#1;data_in = testData5[8663];
@(posedge clk);
#1;data_in = testData5[8664];
@(posedge clk);
#1;data_in = testData5[8665];
@(posedge clk);
#1;data_in = testData5[8666];
@(posedge clk);
#1;data_in = testData5[8667];
@(posedge clk);
#1;data_in = testData5[8668];
@(posedge clk);
#1;data_in = testData5[8669];
@(posedge clk);
#1;data_in = testData5[8670];
@(posedge clk);
#1;data_in = testData5[8671];
@(posedge clk);
#1;data_in = testData5[8672];
@(posedge clk);
#1;data_in = testData5[8673];
@(posedge clk);
#1;data_in = testData5[8674];
@(posedge clk);
#1;data_in = testData5[8675];
@(posedge clk);
#1;data_in = testData5[8676];
@(posedge clk);
#1;data_in = testData5[8677];
@(posedge clk);
#1;data_in = testData5[8678];
@(posedge clk);
#1;data_in = testData5[8679];
@(posedge clk);
#1;data_in = testData5[8680];
@(posedge clk);
#1;data_in = testData5[8681];
@(posedge clk);
#1;data_in = testData5[8682];
@(posedge clk);
#1;data_in = testData5[8683];
@(posedge clk);
#1;data_in = testData5[8684];
@(posedge clk);
#1;data_in = testData5[8685];
@(posedge clk);
#1;data_in = testData5[8686];
@(posedge clk);
#1;data_in = testData5[8687];
@(posedge clk);
#1;data_in = testData5[8688];
@(posedge clk);
#1;data_in = testData5[8689];
@(posedge clk);
#1;data_in = testData5[8690];
@(posedge clk);
#1;data_in = testData5[8691];
@(posedge clk);
#1;data_in = testData5[8692];
@(posedge clk);
#1;data_in = testData5[8693];
@(posedge clk);
#1;data_in = testData5[8694];
@(posedge clk);
#1;data_in = testData5[8695];
@(posedge clk);
#1;data_in = testData5[8696];
@(posedge clk);
#1;data_in = testData5[8697];
@(posedge clk);
#1;data_in = testData5[8698];
@(posedge clk);
#1;data_in = testData5[8699];
@(posedge clk);
#1;data_in = testData5[8700];
@(posedge clk);
#1;data_in = testData5[8701];
@(posedge clk);
#1;data_in = testData5[8702];
@(posedge clk);
#1;data_in = testData5[8703];
@(posedge clk);
#1;data_in = testData5[8704];
@(posedge clk);
#1;data_in = testData5[8705];
@(posedge clk);
#1;data_in = testData5[8706];
@(posedge clk);
#1;data_in = testData5[8707];
@(posedge clk);
#1;data_in = testData5[8708];
@(posedge clk);
#1;data_in = testData5[8709];
@(posedge clk);
#1;data_in = testData5[8710];
@(posedge clk);
#1;data_in = testData5[8711];
@(posedge clk);
#1;data_in = testData5[8712];
@(posedge clk);
#1;data_in = testData5[8713];
@(posedge clk);
#1;data_in = testData5[8714];
@(posedge clk);
#1;data_in = testData5[8715];
@(posedge clk);
#1;data_in = testData5[8716];
@(posedge clk);
#1;data_in = testData5[8717];
@(posedge clk);
#1;data_in = testData5[8718];
@(posedge clk);
#1;data_in = testData5[8719];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[8720]; 
@(posedge clk);
#1;data_in = testData5[8721];
@(posedge clk);
#1;data_in = testData5[8722];
@(posedge clk);
#1;data_in = testData5[8723];
@(posedge clk);
#1;data_in = testData5[8724];
@(posedge clk);
#1;data_in = testData5[8725];
@(posedge clk);
#1;data_in = testData5[8726];
@(posedge clk);
#1;data_in = testData5[8727];
@(posedge clk);
#1;data_in = testData5[8728];
@(posedge clk);
#1;data_in = testData5[8729];
@(posedge clk);
#1;data_in = testData5[8730];
@(posedge clk);
#1;data_in = testData5[8731];
@(posedge clk);
#1;data_in = testData5[8732];
@(posedge clk);
#1;data_in = testData5[8733];
@(posedge clk);
#1;data_in = testData5[8734];
@(posedge clk);
#1;data_in = testData5[8735];
@(posedge clk);
#1;data_in = testData5[8736];
@(posedge clk);
#1;data_in = testData5[8737];
@(posedge clk);
#1;data_in = testData5[8738];
@(posedge clk);
#1;data_in = testData5[8739];
@(posedge clk);
#1;data_in = testData5[8740];
@(posedge clk);
#1;data_in = testData5[8741];
@(posedge clk);
#1;data_in = testData5[8742];
@(posedge clk);
#1;data_in = testData5[8743];
@(posedge clk);
#1;data_in = testData5[8744];
@(posedge clk);
#1;data_in = testData5[8745];
@(posedge clk);
#1;data_in = testData5[8746];
@(posedge clk);
#1;data_in = testData5[8747];
@(posedge clk);
#1;data_in = testData5[8748];
@(posedge clk);
#1;data_in = testData5[8749];
@(posedge clk);
#1;data_in = testData5[8750];
@(posedge clk);
#1;data_in = testData5[8751];
@(posedge clk);
#1;data_in = testData5[8752];
@(posedge clk);
#1;data_in = testData5[8753];
@(posedge clk);
#1;data_in = testData5[8754];
@(posedge clk);
#1;data_in = testData5[8755];
@(posedge clk);
#1;data_in = testData5[8756];
@(posedge clk);
#1;data_in = testData5[8757];
@(posedge clk);
#1;data_in = testData5[8758];
@(posedge clk);
#1;data_in = testData5[8759];
@(posedge clk);
#1;data_in = testData5[8760];
@(posedge clk);
#1;data_in = testData5[8761];
@(posedge clk);
#1;data_in = testData5[8762];
@(posedge clk);
#1;data_in = testData5[8763];
@(posedge clk);
#1;data_in = testData5[8764];
@(posedge clk);
#1;data_in = testData5[8765];
@(posedge clk);
#1;data_in = testData5[8766];
@(posedge clk);
#1;data_in = testData5[8767];
@(posedge clk);
#1;data_in = testData5[8768];
@(posedge clk);
#1;data_in = testData5[8769];
@(posedge clk);
#1;data_in = testData5[8770];
@(posedge clk);
#1;data_in = testData5[8771];
@(posedge clk);
#1;data_in = testData5[8772];
@(posedge clk);
#1;data_in = testData5[8773];
@(posedge clk);
#1;data_in = testData5[8774];
@(posedge clk);
#1;data_in = testData5[8775];
@(posedge clk);
#1;data_in = testData5[8776];
@(posedge clk);
#1;data_in = testData5[8777];
@(posedge clk);
#1;data_in = testData5[8778];
@(posedge clk);
#1;data_in = testData5[8779];
@(posedge clk);
#1;data_in = testData5[8780];
@(posedge clk);
#1;data_in = testData5[8781];
@(posedge clk);
#1;data_in = testData5[8782];
@(posedge clk);
#1;data_in = testData5[8783];
@(posedge clk);
#1;data_in = testData5[8784];
@(posedge clk);
#1;data_in = testData5[8785];
@(posedge clk);
#1;data_in = testData5[8786];
@(posedge clk);
#1;data_in = testData5[8787];
@(posedge clk);
#1;data_in = testData5[8788];
@(posedge clk);
#1;data_in = testData5[8789];
@(posedge clk);
#1;data_in = testData5[8790];
@(posedge clk);
#1;data_in = testData5[8791];
@(posedge clk);
#1;data_in = testData5[8792];
@(posedge clk);
#1;data_in = testData5[8793];
@(posedge clk);
#1;data_in = testData5[8794];
@(posedge clk);
#1;data_in = testData5[8795];
@(posedge clk);
#1;data_in = testData5[8796];
@(posedge clk);
#1;data_in = testData5[8797];
@(posedge clk);
#1;data_in = testData5[8798];
@(posedge clk);
#1;data_in = testData5[8799];
@(posedge clk);
#1;data_in = testData5[8800];
@(posedge clk);
#1;data_in = testData5[8801];
@(posedge clk);
#1;data_in = testData5[8802];
@(posedge clk);
#1;data_in = testData5[8803];
@(posedge clk);
#1;data_in = testData5[8804];
@(posedge clk);
#1;data_in = testData5[8805];
@(posedge clk);
#1;data_in = testData5[8806];
@(posedge clk);
#1;data_in = testData5[8807];
@(posedge clk);
#1;data_in = testData5[8808];
@(posedge clk);
#1;data_in = testData5[8809];
@(posedge clk);
#1;data_in = testData5[8810];
@(posedge clk);
#1;data_in = testData5[8811];
@(posedge clk);
#1;data_in = testData5[8812];
@(posedge clk);
#1;data_in = testData5[8813];
@(posedge clk);
#1;data_in = testData5[8814];
@(posedge clk);
#1;data_in = testData5[8815];
@(posedge clk);
#1;data_in = testData5[8816];
@(posedge clk);
#1;data_in = testData5[8817];
@(posedge clk);
#1;data_in = testData5[8818];
@(posedge clk);
#1;data_in = testData5[8819];
@(posedge clk);
#1;data_in = testData5[8820];
@(posedge clk);
#1;data_in = testData5[8821];
@(posedge clk);
#1;data_in = testData5[8822];
@(posedge clk);
#1;data_in = testData5[8823];
@(posedge clk);
#1;data_in = testData5[8824];
@(posedge clk);
#1;data_in = testData5[8825];
@(posedge clk);
#1;data_in = testData5[8826];
@(posedge clk);
#1;data_in = testData5[8827];
@(posedge clk);
#1;data_in = testData5[8828];
@(posedge clk);
#1;data_in = testData5[8829];
@(posedge clk);
#1;data_in = testData5[8830];
@(posedge clk);
#1;data_in = testData5[8831];
@(posedge clk);
#1;data_in = testData5[8832];
@(posedge clk);
#1;data_in = testData5[8833];
@(posedge clk);
#1;data_in = testData5[8834];
@(posedge clk);
#1;data_in = testData5[8835];
@(posedge clk);
#1;data_in = testData5[8836];
@(posedge clk);
#1;data_in = testData5[8837];
@(posedge clk);
#1;data_in = testData5[8838];
@(posedge clk);
#1;data_in = testData5[8839];
@(posedge clk);
#1;data_in = testData5[8840];
@(posedge clk);
#1;data_in = testData5[8841];
@(posedge clk);
#1;data_in = testData5[8842];
@(posedge clk);
#1;data_in = testData5[8843];
@(posedge clk);
#1;data_in = testData5[8844];
@(posedge clk);
#1;data_in = testData5[8845];
@(posedge clk);
#1;data_in = testData5[8846];
@(posedge clk);
#1;data_in = testData5[8847];
@(posedge clk);
#1;data_in = testData5[8848];
@(posedge clk);
#1;data_in = testData5[8849];
@(posedge clk);
#1;data_in = testData5[8850];
@(posedge clk);
#1;data_in = testData5[8851];
@(posedge clk);
#1;data_in = testData5[8852];
@(posedge clk);
#1;data_in = testData5[8853];
@(posedge clk);
#1;data_in = testData5[8854];
@(posedge clk);
#1;data_in = testData5[8855];
@(posedge clk);
#1;data_in = testData5[8856];
@(posedge clk);
#1;data_in = testData5[8857];
@(posedge clk);
#1;data_in = testData5[8858];
@(posedge clk);
#1;data_in = testData5[8859];
@(posedge clk);
#1;data_in = testData5[8860];
@(posedge clk);
#1;data_in = testData5[8861];
@(posedge clk);
#1;data_in = testData5[8862];
@(posedge clk);
#1;data_in = testData5[8863];
@(posedge clk);
#1;data_in = testData5[8864];
@(posedge clk);
#1;data_in = testData5[8865];
@(posedge clk);
#1;data_in = testData5[8866];
@(posedge clk);
#1;data_in = testData5[8867];
@(posedge clk);
#1;data_in = testData5[8868];
@(posedge clk);
#1;data_in = testData5[8869];
@(posedge clk);
#1;data_in = testData5[8870];
@(posedge clk);
#1;data_in = testData5[8871];
@(posedge clk);
#1;data_in = testData5[8872];
@(posedge clk);
#1;data_in = testData5[8873];
@(posedge clk);
#1;data_in = testData5[8874];
@(posedge clk);
#1;data_in = testData5[8875];
@(posedge clk);
#1;data_in = testData5[8876];
@(posedge clk);
#1;data_in = testData5[8877];
@(posedge clk);
#1;data_in = testData5[8878];
@(posedge clk);
#1;data_in = testData5[8879];
@(posedge clk);
#1;data_in = testData5[8880];
@(posedge clk);
#1;data_in = testData5[8881];
@(posedge clk);
#1;data_in = testData5[8882];
@(posedge clk);
#1;data_in = testData5[8883];
@(posedge clk);
#1;data_in = testData5[8884];
@(posedge clk);
#1;data_in = testData5[8885];
@(posedge clk);
#1;data_in = testData5[8886];
@(posedge clk);
#1;data_in = testData5[8887];
@(posedge clk);
#1;data_in = testData5[8888];
@(posedge clk);
#1;data_in = testData5[8889];
@(posedge clk);
#1;data_in = testData5[8890];
@(posedge clk);
#1;data_in = testData5[8891];
@(posedge clk);
#1;data_in = testData5[8892];
@(posedge clk);
#1;data_in = testData5[8893];
@(posedge clk);
#1;data_in = testData5[8894];
@(posedge clk);
#1;data_in = testData5[8895];
@(posedge clk);
#1;data_in = testData5[8896];
@(posedge clk);
#1;data_in = testData5[8897];
@(posedge clk);
#1;data_in = testData5[8898];
@(posedge clk);
#1;data_in = testData5[8899];
@(posedge clk);
#1;data_in = testData5[8900];
@(posedge clk);
#1;data_in = testData5[8901];
@(posedge clk);
#1;data_in = testData5[8902];
@(posedge clk);
#1;data_in = testData5[8903];
@(posedge clk);
#1;data_in = testData5[8904];
@(posedge clk);
#1;data_in = testData5[8905];
@(posedge clk);
#1;data_in = testData5[8906];
@(posedge clk);
#1;data_in = testData5[8907];
@(posedge clk);
#1;data_in = testData5[8908];
@(posedge clk);
#1;data_in = testData5[8909];
@(posedge clk);
#1;data_in = testData5[8910];
@(posedge clk);
#1;data_in = testData5[8911];
@(posedge clk);
#1;data_in = testData5[8912];
@(posedge clk);
#1;data_in = testData5[8913];
@(posedge clk);
#1;data_in = testData5[8914];
@(posedge clk);
#1;data_in = testData5[8915];
@(posedge clk);
#1;data_in = testData5[8916];
@(posedge clk);
#1;data_in = testData5[8917];
@(posedge clk);
#1;data_in = testData5[8918];
@(posedge clk);
#1;data_in = testData5[8919];
@(posedge clk);
#1;data_in = testData5[8920];
@(posedge clk);
#1;data_in = testData5[8921];
@(posedge clk);
#1;data_in = testData5[8922];
@(posedge clk);
#1;data_in = testData5[8923];
@(posedge clk);
#1;data_in = testData5[8924];
@(posedge clk);
#1;data_in = testData5[8925];
@(posedge clk);
#1;data_in = testData5[8926];
@(posedge clk);
#1;data_in = testData5[8927];
@(posedge clk);
#1;data_in = testData5[8928];
@(posedge clk);
#1;data_in = testData5[8929];
@(posedge clk);
#1;data_in = testData5[8930];
@(posedge clk);
#1;data_in = testData5[8931];
@(posedge clk);
#1;data_in = testData5[8932];
@(posedge clk);
#1;data_in = testData5[8933];
@(posedge clk);
#1;data_in = testData5[8934];
@(posedge clk);
#1;data_in = testData5[8935];
@(posedge clk);
#1;data_in = testData5[8936];
@(posedge clk);
#1;data_in = testData5[8937];
@(posedge clk);
#1;data_in = testData5[8938];
@(posedge clk);
#1;data_in = testData5[8939];
@(posedge clk);
#1;data_in = testData5[8940];
@(posedge clk);
#1;data_in = testData5[8941];
@(posedge clk);
#1;data_in = testData5[8942];
@(posedge clk);
#1;data_in = testData5[8943];
@(posedge clk);
#1;data_in = testData5[8944];
@(posedge clk);
#1;data_in = testData5[8945];
@(posedge clk);
#1;data_in = testData5[8946];
@(posedge clk);
#1;data_in = testData5[8947];
@(posedge clk);
#1;data_in = testData5[8948];
@(posedge clk);
#1;data_in = testData5[8949];
@(posedge clk);
#1;data_in = testData5[8950];
@(posedge clk);
#1;data_in = testData5[8951];
@(posedge clk);
#1;data_in = testData5[8952];
@(posedge clk);
#1;data_in = testData5[8953];
@(posedge clk);
#1;data_in = testData5[8954];
@(posedge clk);
#1;data_in = testData5[8955];
@(posedge clk);
#1;data_in = testData5[8956];
@(posedge clk);
#1;data_in = testData5[8957];
@(posedge clk);
#1;data_in = testData5[8958];
@(posedge clk);
#1;data_in = testData5[8959];
@(posedge clk);
#1;data_in = testData5[8960];
@(posedge clk);
#1;data_in = testData5[8961];
@(posedge clk);
#1;data_in = testData5[8962];
@(posedge clk);
#1;data_in = testData5[8963];
@(posedge clk);
#1;data_in = testData5[8964];
@(posedge clk);
#1;data_in = testData5[8965];
@(posedge clk);
#1;data_in = testData5[8966];
@(posedge clk);
#1;data_in = testData5[8967];
@(posedge clk);
#1;data_in = testData5[8968];
@(posedge clk);
#1;data_in = testData5[8969];
@(posedge clk);
#1;data_in = testData5[8970];
@(posedge clk);
#1;data_in = testData5[8971];
@(posedge clk);
#1;data_in = testData5[8972];
@(posedge clk);
#1;data_in = testData5[8973];
@(posedge clk);
#1;data_in = testData5[8974];
@(posedge clk);
#1;data_in = testData5[8975];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[8976]; 
@(posedge clk);
#1;data_in = testData5[8977];
@(posedge clk);
#1;data_in = testData5[8978];
@(posedge clk);
#1;data_in = testData5[8979];
@(posedge clk);
#1;data_in = testData5[8980];
@(posedge clk);
#1;data_in = testData5[8981];
@(posedge clk);
#1;data_in = testData5[8982];
@(posedge clk);
#1;data_in = testData5[8983];
@(posedge clk);
#1;data_in = testData5[8984];
@(posedge clk);
#1;data_in = testData5[8985];
@(posedge clk);
#1;data_in = testData5[8986];
@(posedge clk);
#1;data_in = testData5[8987];
@(posedge clk);
#1;data_in = testData5[8988];
@(posedge clk);
#1;data_in = testData5[8989];
@(posedge clk);
#1;data_in = testData5[8990];
@(posedge clk);
#1;data_in = testData5[8991];
@(posedge clk);
#1;data_in = testData5[8992];
@(posedge clk);
#1;data_in = testData5[8993];
@(posedge clk);
#1;data_in = testData5[8994];
@(posedge clk);
#1;data_in = testData5[8995];
@(posedge clk);
#1;data_in = testData5[8996];
@(posedge clk);
#1;data_in = testData5[8997];
@(posedge clk);
#1;data_in = testData5[8998];
@(posedge clk);
#1;data_in = testData5[8999];
@(posedge clk);
#1;data_in = testData5[9000];
@(posedge clk);
#1;data_in = testData5[9001];
@(posedge clk);
#1;data_in = testData5[9002];
@(posedge clk);
#1;data_in = testData5[9003];
@(posedge clk);
#1;data_in = testData5[9004];
@(posedge clk);
#1;data_in = testData5[9005];
@(posedge clk);
#1;data_in = testData5[9006];
@(posedge clk);
#1;data_in = testData5[9007];
@(posedge clk);
#1;data_in = testData5[9008];
@(posedge clk);
#1;data_in = testData5[9009];
@(posedge clk);
#1;data_in = testData5[9010];
@(posedge clk);
#1;data_in = testData5[9011];
@(posedge clk);
#1;data_in = testData5[9012];
@(posedge clk);
#1;data_in = testData5[9013];
@(posedge clk);
#1;data_in = testData5[9014];
@(posedge clk);
#1;data_in = testData5[9015];
@(posedge clk);
#1;data_in = testData5[9016];
@(posedge clk);
#1;data_in = testData5[9017];
@(posedge clk);
#1;data_in = testData5[9018];
@(posedge clk);
#1;data_in = testData5[9019];
@(posedge clk);
#1;data_in = testData5[9020];
@(posedge clk);
#1;data_in = testData5[9021];
@(posedge clk);
#1;data_in = testData5[9022];
@(posedge clk);
#1;data_in = testData5[9023];
@(posedge clk);
#1;data_in = testData5[9024];
@(posedge clk);
#1;data_in = testData5[9025];
@(posedge clk);
#1;data_in = testData5[9026];
@(posedge clk);
#1;data_in = testData5[9027];
@(posedge clk);
#1;data_in = testData5[9028];
@(posedge clk);
#1;data_in = testData5[9029];
@(posedge clk);
#1;data_in = testData5[9030];
@(posedge clk);
#1;data_in = testData5[9031];
@(posedge clk);
#1;data_in = testData5[9032];
@(posedge clk);
#1;data_in = testData5[9033];
@(posedge clk);
#1;data_in = testData5[9034];
@(posedge clk);
#1;data_in = testData5[9035];
@(posedge clk);
#1;data_in = testData5[9036];
@(posedge clk);
#1;data_in = testData5[9037];
@(posedge clk);
#1;data_in = testData5[9038];
@(posedge clk);
#1;data_in = testData5[9039];
@(posedge clk);
#1;data_in = testData5[9040];
@(posedge clk);
#1;data_in = testData5[9041];
@(posedge clk);
#1;data_in = testData5[9042];
@(posedge clk);
#1;data_in = testData5[9043];
@(posedge clk);
#1;data_in = testData5[9044];
@(posedge clk);
#1;data_in = testData5[9045];
@(posedge clk);
#1;data_in = testData5[9046];
@(posedge clk);
#1;data_in = testData5[9047];
@(posedge clk);
#1;data_in = testData5[9048];
@(posedge clk);
#1;data_in = testData5[9049];
@(posedge clk);
#1;data_in = testData5[9050];
@(posedge clk);
#1;data_in = testData5[9051];
@(posedge clk);
#1;data_in = testData5[9052];
@(posedge clk);
#1;data_in = testData5[9053];
@(posedge clk);
#1;data_in = testData5[9054];
@(posedge clk);
#1;data_in = testData5[9055];
@(posedge clk);
#1;data_in = testData5[9056];
@(posedge clk);
#1;data_in = testData5[9057];
@(posedge clk);
#1;data_in = testData5[9058];
@(posedge clk);
#1;data_in = testData5[9059];
@(posedge clk);
#1;data_in = testData5[9060];
@(posedge clk);
#1;data_in = testData5[9061];
@(posedge clk);
#1;data_in = testData5[9062];
@(posedge clk);
#1;data_in = testData5[9063];
@(posedge clk);
#1;data_in = testData5[9064];
@(posedge clk);
#1;data_in = testData5[9065];
@(posedge clk);
#1;data_in = testData5[9066];
@(posedge clk);
#1;data_in = testData5[9067];
@(posedge clk);
#1;data_in = testData5[9068];
@(posedge clk);
#1;data_in = testData5[9069];
@(posedge clk);
#1;data_in = testData5[9070];
@(posedge clk);
#1;data_in = testData5[9071];
@(posedge clk);
#1;data_in = testData5[9072];
@(posedge clk);
#1;data_in = testData5[9073];
@(posedge clk);
#1;data_in = testData5[9074];
@(posedge clk);
#1;data_in = testData5[9075];
@(posedge clk);
#1;data_in = testData5[9076];
@(posedge clk);
#1;data_in = testData5[9077];
@(posedge clk);
#1;data_in = testData5[9078];
@(posedge clk);
#1;data_in = testData5[9079];
@(posedge clk);
#1;data_in = testData5[9080];
@(posedge clk);
#1;data_in = testData5[9081];
@(posedge clk);
#1;data_in = testData5[9082];
@(posedge clk);
#1;data_in = testData5[9083];
@(posedge clk);
#1;data_in = testData5[9084];
@(posedge clk);
#1;data_in = testData5[9085];
@(posedge clk);
#1;data_in = testData5[9086];
@(posedge clk);
#1;data_in = testData5[9087];
@(posedge clk);
#1;data_in = testData5[9088];
@(posedge clk);
#1;data_in = testData5[9089];
@(posedge clk);
#1;data_in = testData5[9090];
@(posedge clk);
#1;data_in = testData5[9091];
@(posedge clk);
#1;data_in = testData5[9092];
@(posedge clk);
#1;data_in = testData5[9093];
@(posedge clk);
#1;data_in = testData5[9094];
@(posedge clk);
#1;data_in = testData5[9095];
@(posedge clk);
#1;data_in = testData5[9096];
@(posedge clk);
#1;data_in = testData5[9097];
@(posedge clk);
#1;data_in = testData5[9098];
@(posedge clk);
#1;data_in = testData5[9099];
@(posedge clk);
#1;data_in = testData5[9100];
@(posedge clk);
#1;data_in = testData5[9101];
@(posedge clk);
#1;data_in = testData5[9102];
@(posedge clk);
#1;data_in = testData5[9103];
@(posedge clk);
#1;data_in = testData5[9104];
@(posedge clk);
#1;data_in = testData5[9105];
@(posedge clk);
#1;data_in = testData5[9106];
@(posedge clk);
#1;data_in = testData5[9107];
@(posedge clk);
#1;data_in = testData5[9108];
@(posedge clk);
#1;data_in = testData5[9109];
@(posedge clk);
#1;data_in = testData5[9110];
@(posedge clk);
#1;data_in = testData5[9111];
@(posedge clk);
#1;data_in = testData5[9112];
@(posedge clk);
#1;data_in = testData5[9113];
@(posedge clk);
#1;data_in = testData5[9114];
@(posedge clk);
#1;data_in = testData5[9115];
@(posedge clk);
#1;data_in = testData5[9116];
@(posedge clk);
#1;data_in = testData5[9117];
@(posedge clk);
#1;data_in = testData5[9118];
@(posedge clk);
#1;data_in = testData5[9119];
@(posedge clk);
#1;data_in = testData5[9120];
@(posedge clk);
#1;data_in = testData5[9121];
@(posedge clk);
#1;data_in = testData5[9122];
@(posedge clk);
#1;data_in = testData5[9123];
@(posedge clk);
#1;data_in = testData5[9124];
@(posedge clk);
#1;data_in = testData5[9125];
@(posedge clk);
#1;data_in = testData5[9126];
@(posedge clk);
#1;data_in = testData5[9127];
@(posedge clk);
#1;data_in = testData5[9128];
@(posedge clk);
#1;data_in = testData5[9129];
@(posedge clk);
#1;data_in = testData5[9130];
@(posedge clk);
#1;data_in = testData5[9131];
@(posedge clk);
#1;data_in = testData5[9132];
@(posedge clk);
#1;data_in = testData5[9133];
@(posedge clk);
#1;data_in = testData5[9134];
@(posedge clk);
#1;data_in = testData5[9135];
@(posedge clk);
#1;data_in = testData5[9136];
@(posedge clk);
#1;data_in = testData5[9137];
@(posedge clk);
#1;data_in = testData5[9138];
@(posedge clk);
#1;data_in = testData5[9139];
@(posedge clk);
#1;data_in = testData5[9140];
@(posedge clk);
#1;data_in = testData5[9141];
@(posedge clk);
#1;data_in = testData5[9142];
@(posedge clk);
#1;data_in = testData5[9143];
@(posedge clk);
#1;data_in = testData5[9144];
@(posedge clk);
#1;data_in = testData5[9145];
@(posedge clk);
#1;data_in = testData5[9146];
@(posedge clk);
#1;data_in = testData5[9147];
@(posedge clk);
#1;data_in = testData5[9148];
@(posedge clk);
#1;data_in = testData5[9149];
@(posedge clk);
#1;data_in = testData5[9150];
@(posedge clk);
#1;data_in = testData5[9151];
@(posedge clk);
#1;data_in = testData5[9152];
@(posedge clk);
#1;data_in = testData5[9153];
@(posedge clk);
#1;data_in = testData5[9154];
@(posedge clk);
#1;data_in = testData5[9155];
@(posedge clk);
#1;data_in = testData5[9156];
@(posedge clk);
#1;data_in = testData5[9157];
@(posedge clk);
#1;data_in = testData5[9158];
@(posedge clk);
#1;data_in = testData5[9159];
@(posedge clk);
#1;data_in = testData5[9160];
@(posedge clk);
#1;data_in = testData5[9161];
@(posedge clk);
#1;data_in = testData5[9162];
@(posedge clk);
#1;data_in = testData5[9163];
@(posedge clk);
#1;data_in = testData5[9164];
@(posedge clk);
#1;data_in = testData5[9165];
@(posedge clk);
#1;data_in = testData5[9166];
@(posedge clk);
#1;data_in = testData5[9167];
@(posedge clk);
#1;data_in = testData5[9168];
@(posedge clk);
#1;data_in = testData5[9169];
@(posedge clk);
#1;data_in = testData5[9170];
@(posedge clk);
#1;data_in = testData5[9171];
@(posedge clk);
#1;data_in = testData5[9172];
@(posedge clk);
#1;data_in = testData5[9173];
@(posedge clk);
#1;data_in = testData5[9174];
@(posedge clk);
#1;data_in = testData5[9175];
@(posedge clk);
#1;data_in = testData5[9176];
@(posedge clk);
#1;data_in = testData5[9177];
@(posedge clk);
#1;data_in = testData5[9178];
@(posedge clk);
#1;data_in = testData5[9179];
@(posedge clk);
#1;data_in = testData5[9180];
@(posedge clk);
#1;data_in = testData5[9181];
@(posedge clk);
#1;data_in = testData5[9182];
@(posedge clk);
#1;data_in = testData5[9183];
@(posedge clk);
#1;data_in = testData5[9184];
@(posedge clk);
#1;data_in = testData5[9185];
@(posedge clk);
#1;data_in = testData5[9186];
@(posedge clk);
#1;data_in = testData5[9187];
@(posedge clk);
#1;data_in = testData5[9188];
@(posedge clk);
#1;data_in = testData5[9189];
@(posedge clk);
#1;data_in = testData5[9190];
@(posedge clk);
#1;data_in = testData5[9191];
@(posedge clk);
#1;data_in = testData5[9192];
@(posedge clk);
#1;data_in = testData5[9193];
@(posedge clk);
#1;data_in = testData5[9194];
@(posedge clk);
#1;data_in = testData5[9195];
@(posedge clk);
#1;data_in = testData5[9196];
@(posedge clk);
#1;data_in = testData5[9197];
@(posedge clk);
#1;data_in = testData5[9198];
@(posedge clk);
#1;data_in = testData5[9199];
@(posedge clk);
#1;data_in = testData5[9200];
@(posedge clk);
#1;data_in = testData5[9201];
@(posedge clk);
#1;data_in = testData5[9202];
@(posedge clk);
#1;data_in = testData5[9203];
@(posedge clk);
#1;data_in = testData5[9204];
@(posedge clk);
#1;data_in = testData5[9205];
@(posedge clk);
#1;data_in = testData5[9206];
@(posedge clk);
#1;data_in = testData5[9207];
@(posedge clk);
#1;data_in = testData5[9208];
@(posedge clk);
#1;data_in = testData5[9209];
@(posedge clk);
#1;data_in = testData5[9210];
@(posedge clk);
#1;data_in = testData5[9211];
@(posedge clk);
#1;data_in = testData5[9212];
@(posedge clk);
#1;data_in = testData5[9213];
@(posedge clk);
#1;data_in = testData5[9214];
@(posedge clk);
#1;data_in = testData5[9215];
@(posedge clk);
#1;data_in = testData5[9216];
@(posedge clk);
#1;data_in = testData5[9217];
@(posedge clk);
#1;data_in = testData5[9218];
@(posedge clk);
#1;data_in = testData5[9219];
@(posedge clk);
#1;data_in = testData5[9220];
@(posedge clk);
#1;data_in = testData5[9221];
@(posedge clk);
#1;data_in = testData5[9222];
@(posedge clk);
#1;data_in = testData5[9223];
@(posedge clk);
#1;data_in = testData5[9224];
@(posedge clk);
#1;data_in = testData5[9225];
@(posedge clk);
#1;data_in = testData5[9226];
@(posedge clk);
#1;data_in = testData5[9227];
@(posedge clk);
#1;data_in = testData5[9228];
@(posedge clk);
#1;data_in = testData5[9229];
@(posedge clk);
#1;data_in = testData5[9230];
@(posedge clk);
#1;data_in = testData5[9231];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[9232]; 
@(posedge clk);
#1;data_in = testData5[9233];
@(posedge clk);
#1;data_in = testData5[9234];
@(posedge clk);
#1;data_in = testData5[9235];
@(posedge clk);
#1;data_in = testData5[9236];
@(posedge clk);
#1;data_in = testData5[9237];
@(posedge clk);
#1;data_in = testData5[9238];
@(posedge clk);
#1;data_in = testData5[9239];
@(posedge clk);
#1;data_in = testData5[9240];
@(posedge clk);
#1;data_in = testData5[9241];
@(posedge clk);
#1;data_in = testData5[9242];
@(posedge clk);
#1;data_in = testData5[9243];
@(posedge clk);
#1;data_in = testData5[9244];
@(posedge clk);
#1;data_in = testData5[9245];
@(posedge clk);
#1;data_in = testData5[9246];
@(posedge clk);
#1;data_in = testData5[9247];
@(posedge clk);
#1;data_in = testData5[9248];
@(posedge clk);
#1;data_in = testData5[9249];
@(posedge clk);
#1;data_in = testData5[9250];
@(posedge clk);
#1;data_in = testData5[9251];
@(posedge clk);
#1;data_in = testData5[9252];
@(posedge clk);
#1;data_in = testData5[9253];
@(posedge clk);
#1;data_in = testData5[9254];
@(posedge clk);
#1;data_in = testData5[9255];
@(posedge clk);
#1;data_in = testData5[9256];
@(posedge clk);
#1;data_in = testData5[9257];
@(posedge clk);
#1;data_in = testData5[9258];
@(posedge clk);
#1;data_in = testData5[9259];
@(posedge clk);
#1;data_in = testData5[9260];
@(posedge clk);
#1;data_in = testData5[9261];
@(posedge clk);
#1;data_in = testData5[9262];
@(posedge clk);
#1;data_in = testData5[9263];
@(posedge clk);
#1;data_in = testData5[9264];
@(posedge clk);
#1;data_in = testData5[9265];
@(posedge clk);
#1;data_in = testData5[9266];
@(posedge clk);
#1;data_in = testData5[9267];
@(posedge clk);
#1;data_in = testData5[9268];
@(posedge clk);
#1;data_in = testData5[9269];
@(posedge clk);
#1;data_in = testData5[9270];
@(posedge clk);
#1;data_in = testData5[9271];
@(posedge clk);
#1;data_in = testData5[9272];
@(posedge clk);
#1;data_in = testData5[9273];
@(posedge clk);
#1;data_in = testData5[9274];
@(posedge clk);
#1;data_in = testData5[9275];
@(posedge clk);
#1;data_in = testData5[9276];
@(posedge clk);
#1;data_in = testData5[9277];
@(posedge clk);
#1;data_in = testData5[9278];
@(posedge clk);
#1;data_in = testData5[9279];
@(posedge clk);
#1;data_in = testData5[9280];
@(posedge clk);
#1;data_in = testData5[9281];
@(posedge clk);
#1;data_in = testData5[9282];
@(posedge clk);
#1;data_in = testData5[9283];
@(posedge clk);
#1;data_in = testData5[9284];
@(posedge clk);
#1;data_in = testData5[9285];
@(posedge clk);
#1;data_in = testData5[9286];
@(posedge clk);
#1;data_in = testData5[9287];
@(posedge clk);
#1;data_in = testData5[9288];
@(posedge clk);
#1;data_in = testData5[9289];
@(posedge clk);
#1;data_in = testData5[9290];
@(posedge clk);
#1;data_in = testData5[9291];
@(posedge clk);
#1;data_in = testData5[9292];
@(posedge clk);
#1;data_in = testData5[9293];
@(posedge clk);
#1;data_in = testData5[9294];
@(posedge clk);
#1;data_in = testData5[9295];
@(posedge clk);
#1;data_in = testData5[9296];
@(posedge clk);
#1;data_in = testData5[9297];
@(posedge clk);
#1;data_in = testData5[9298];
@(posedge clk);
#1;data_in = testData5[9299];
@(posedge clk);
#1;data_in = testData5[9300];
@(posedge clk);
#1;data_in = testData5[9301];
@(posedge clk);
#1;data_in = testData5[9302];
@(posedge clk);
#1;data_in = testData5[9303];
@(posedge clk);
#1;data_in = testData5[9304];
@(posedge clk);
#1;data_in = testData5[9305];
@(posedge clk);
#1;data_in = testData5[9306];
@(posedge clk);
#1;data_in = testData5[9307];
@(posedge clk);
#1;data_in = testData5[9308];
@(posedge clk);
#1;data_in = testData5[9309];
@(posedge clk);
#1;data_in = testData5[9310];
@(posedge clk);
#1;data_in = testData5[9311];
@(posedge clk);
#1;data_in = testData5[9312];
@(posedge clk);
#1;data_in = testData5[9313];
@(posedge clk);
#1;data_in = testData5[9314];
@(posedge clk);
#1;data_in = testData5[9315];
@(posedge clk);
#1;data_in = testData5[9316];
@(posedge clk);
#1;data_in = testData5[9317];
@(posedge clk);
#1;data_in = testData5[9318];
@(posedge clk);
#1;data_in = testData5[9319];
@(posedge clk);
#1;data_in = testData5[9320];
@(posedge clk);
#1;data_in = testData5[9321];
@(posedge clk);
#1;data_in = testData5[9322];
@(posedge clk);
#1;data_in = testData5[9323];
@(posedge clk);
#1;data_in = testData5[9324];
@(posedge clk);
#1;data_in = testData5[9325];
@(posedge clk);
#1;data_in = testData5[9326];
@(posedge clk);
#1;data_in = testData5[9327];
@(posedge clk);
#1;data_in = testData5[9328];
@(posedge clk);
#1;data_in = testData5[9329];
@(posedge clk);
#1;data_in = testData5[9330];
@(posedge clk);
#1;data_in = testData5[9331];
@(posedge clk);
#1;data_in = testData5[9332];
@(posedge clk);
#1;data_in = testData5[9333];
@(posedge clk);
#1;data_in = testData5[9334];
@(posedge clk);
#1;data_in = testData5[9335];
@(posedge clk);
#1;data_in = testData5[9336];
@(posedge clk);
#1;data_in = testData5[9337];
@(posedge clk);
#1;data_in = testData5[9338];
@(posedge clk);
#1;data_in = testData5[9339];
@(posedge clk);
#1;data_in = testData5[9340];
@(posedge clk);
#1;data_in = testData5[9341];
@(posedge clk);
#1;data_in = testData5[9342];
@(posedge clk);
#1;data_in = testData5[9343];
@(posedge clk);
#1;data_in = testData5[9344];
@(posedge clk);
#1;data_in = testData5[9345];
@(posedge clk);
#1;data_in = testData5[9346];
@(posedge clk);
#1;data_in = testData5[9347];
@(posedge clk);
#1;data_in = testData5[9348];
@(posedge clk);
#1;data_in = testData5[9349];
@(posedge clk);
#1;data_in = testData5[9350];
@(posedge clk);
#1;data_in = testData5[9351];
@(posedge clk);
#1;data_in = testData5[9352];
@(posedge clk);
#1;data_in = testData5[9353];
@(posedge clk);
#1;data_in = testData5[9354];
@(posedge clk);
#1;data_in = testData5[9355];
@(posedge clk);
#1;data_in = testData5[9356];
@(posedge clk);
#1;data_in = testData5[9357];
@(posedge clk);
#1;data_in = testData5[9358];
@(posedge clk);
#1;data_in = testData5[9359];
@(posedge clk);
#1;data_in = testData5[9360];
@(posedge clk);
#1;data_in = testData5[9361];
@(posedge clk);
#1;data_in = testData5[9362];
@(posedge clk);
#1;data_in = testData5[9363];
@(posedge clk);
#1;data_in = testData5[9364];
@(posedge clk);
#1;data_in = testData5[9365];
@(posedge clk);
#1;data_in = testData5[9366];
@(posedge clk);
#1;data_in = testData5[9367];
@(posedge clk);
#1;data_in = testData5[9368];
@(posedge clk);
#1;data_in = testData5[9369];
@(posedge clk);
#1;data_in = testData5[9370];
@(posedge clk);
#1;data_in = testData5[9371];
@(posedge clk);
#1;data_in = testData5[9372];
@(posedge clk);
#1;data_in = testData5[9373];
@(posedge clk);
#1;data_in = testData5[9374];
@(posedge clk);
#1;data_in = testData5[9375];
@(posedge clk);
#1;data_in = testData5[9376];
@(posedge clk);
#1;data_in = testData5[9377];
@(posedge clk);
#1;data_in = testData5[9378];
@(posedge clk);
#1;data_in = testData5[9379];
@(posedge clk);
#1;data_in = testData5[9380];
@(posedge clk);
#1;data_in = testData5[9381];
@(posedge clk);
#1;data_in = testData5[9382];
@(posedge clk);
#1;data_in = testData5[9383];
@(posedge clk);
#1;data_in = testData5[9384];
@(posedge clk);
#1;data_in = testData5[9385];
@(posedge clk);
#1;data_in = testData5[9386];
@(posedge clk);
#1;data_in = testData5[9387];
@(posedge clk);
#1;data_in = testData5[9388];
@(posedge clk);
#1;data_in = testData5[9389];
@(posedge clk);
#1;data_in = testData5[9390];
@(posedge clk);
#1;data_in = testData5[9391];
@(posedge clk);
#1;data_in = testData5[9392];
@(posedge clk);
#1;data_in = testData5[9393];
@(posedge clk);
#1;data_in = testData5[9394];
@(posedge clk);
#1;data_in = testData5[9395];
@(posedge clk);
#1;data_in = testData5[9396];
@(posedge clk);
#1;data_in = testData5[9397];
@(posedge clk);
#1;data_in = testData5[9398];
@(posedge clk);
#1;data_in = testData5[9399];
@(posedge clk);
#1;data_in = testData5[9400];
@(posedge clk);
#1;data_in = testData5[9401];
@(posedge clk);
#1;data_in = testData5[9402];
@(posedge clk);
#1;data_in = testData5[9403];
@(posedge clk);
#1;data_in = testData5[9404];
@(posedge clk);
#1;data_in = testData5[9405];
@(posedge clk);
#1;data_in = testData5[9406];
@(posedge clk);
#1;data_in = testData5[9407];
@(posedge clk);
#1;data_in = testData5[9408];
@(posedge clk);
#1;data_in = testData5[9409];
@(posedge clk);
#1;data_in = testData5[9410];
@(posedge clk);
#1;data_in = testData5[9411];
@(posedge clk);
#1;data_in = testData5[9412];
@(posedge clk);
#1;data_in = testData5[9413];
@(posedge clk);
#1;data_in = testData5[9414];
@(posedge clk);
#1;data_in = testData5[9415];
@(posedge clk);
#1;data_in = testData5[9416];
@(posedge clk);
#1;data_in = testData5[9417];
@(posedge clk);
#1;data_in = testData5[9418];
@(posedge clk);
#1;data_in = testData5[9419];
@(posedge clk);
#1;data_in = testData5[9420];
@(posedge clk);
#1;data_in = testData5[9421];
@(posedge clk);
#1;data_in = testData5[9422];
@(posedge clk);
#1;data_in = testData5[9423];
@(posedge clk);
#1;data_in = testData5[9424];
@(posedge clk);
#1;data_in = testData5[9425];
@(posedge clk);
#1;data_in = testData5[9426];
@(posedge clk);
#1;data_in = testData5[9427];
@(posedge clk);
#1;data_in = testData5[9428];
@(posedge clk);
#1;data_in = testData5[9429];
@(posedge clk);
#1;data_in = testData5[9430];
@(posedge clk);
#1;data_in = testData5[9431];
@(posedge clk);
#1;data_in = testData5[9432];
@(posedge clk);
#1;data_in = testData5[9433];
@(posedge clk);
#1;data_in = testData5[9434];
@(posedge clk);
#1;data_in = testData5[9435];
@(posedge clk);
#1;data_in = testData5[9436];
@(posedge clk);
#1;data_in = testData5[9437];
@(posedge clk);
#1;data_in = testData5[9438];
@(posedge clk);
#1;data_in = testData5[9439];
@(posedge clk);
#1;data_in = testData5[9440];
@(posedge clk);
#1;data_in = testData5[9441];
@(posedge clk);
#1;data_in = testData5[9442];
@(posedge clk);
#1;data_in = testData5[9443];
@(posedge clk);
#1;data_in = testData5[9444];
@(posedge clk);
#1;data_in = testData5[9445];
@(posedge clk);
#1;data_in = testData5[9446];
@(posedge clk);
#1;data_in = testData5[9447];
@(posedge clk);
#1;data_in = testData5[9448];
@(posedge clk);
#1;data_in = testData5[9449];
@(posedge clk);
#1;data_in = testData5[9450];
@(posedge clk);
#1;data_in = testData5[9451];
@(posedge clk);
#1;data_in = testData5[9452];
@(posedge clk);
#1;data_in = testData5[9453];
@(posedge clk);
#1;data_in = testData5[9454];
@(posedge clk);
#1;data_in = testData5[9455];
@(posedge clk);
#1;data_in = testData5[9456];
@(posedge clk);
#1;data_in = testData5[9457];
@(posedge clk);
#1;data_in = testData5[9458];
@(posedge clk);
#1;data_in = testData5[9459];
@(posedge clk);
#1;data_in = testData5[9460];
@(posedge clk);
#1;data_in = testData5[9461];
@(posedge clk);
#1;data_in = testData5[9462];
@(posedge clk);
#1;data_in = testData5[9463];
@(posedge clk);
#1;data_in = testData5[9464];
@(posedge clk);
#1;data_in = testData5[9465];
@(posedge clk);
#1;data_in = testData5[9466];
@(posedge clk);
#1;data_in = testData5[9467];
@(posedge clk);
#1;data_in = testData5[9468];
@(posedge clk);
#1;data_in = testData5[9469];
@(posedge clk);
#1;data_in = testData5[9470];
@(posedge clk);
#1;data_in = testData5[9471];
@(posedge clk);
#1;data_in = testData5[9472];
@(posedge clk);
#1;data_in = testData5[9473];
@(posedge clk);
#1;data_in = testData5[9474];
@(posedge clk);
#1;data_in = testData5[9475];
@(posedge clk);
#1;data_in = testData5[9476];
@(posedge clk);
#1;data_in = testData5[9477];
@(posedge clk);
#1;data_in = testData5[9478];
@(posedge clk);
#1;data_in = testData5[9479];
@(posedge clk);
#1;data_in = testData5[9480];
@(posedge clk);
#1;data_in = testData5[9481];
@(posedge clk);
#1;data_in = testData5[9482];
@(posedge clk);
#1;data_in = testData5[9483];
@(posedge clk);
#1;data_in = testData5[9484];
@(posedge clk);
#1;data_in = testData5[9485];
@(posedge clk);
#1;data_in = testData5[9486];
@(posedge clk);
#1;data_in = testData5[9487];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[9488]; 
@(posedge clk);
#1;data_in = testData5[9489];
@(posedge clk);
#1;data_in = testData5[9490];
@(posedge clk);
#1;data_in = testData5[9491];
@(posedge clk);
#1;data_in = testData5[9492];
@(posedge clk);
#1;data_in = testData5[9493];
@(posedge clk);
#1;data_in = testData5[9494];
@(posedge clk);
#1;data_in = testData5[9495];
@(posedge clk);
#1;data_in = testData5[9496];
@(posedge clk);
#1;data_in = testData5[9497];
@(posedge clk);
#1;data_in = testData5[9498];
@(posedge clk);
#1;data_in = testData5[9499];
@(posedge clk);
#1;data_in = testData5[9500];
@(posedge clk);
#1;data_in = testData5[9501];
@(posedge clk);
#1;data_in = testData5[9502];
@(posedge clk);
#1;data_in = testData5[9503];
@(posedge clk);
#1;data_in = testData5[9504];
@(posedge clk);
#1;data_in = testData5[9505];
@(posedge clk);
#1;data_in = testData5[9506];
@(posedge clk);
#1;data_in = testData5[9507];
@(posedge clk);
#1;data_in = testData5[9508];
@(posedge clk);
#1;data_in = testData5[9509];
@(posedge clk);
#1;data_in = testData5[9510];
@(posedge clk);
#1;data_in = testData5[9511];
@(posedge clk);
#1;data_in = testData5[9512];
@(posedge clk);
#1;data_in = testData5[9513];
@(posedge clk);
#1;data_in = testData5[9514];
@(posedge clk);
#1;data_in = testData5[9515];
@(posedge clk);
#1;data_in = testData5[9516];
@(posedge clk);
#1;data_in = testData5[9517];
@(posedge clk);
#1;data_in = testData5[9518];
@(posedge clk);
#1;data_in = testData5[9519];
@(posedge clk);
#1;data_in = testData5[9520];
@(posedge clk);
#1;data_in = testData5[9521];
@(posedge clk);
#1;data_in = testData5[9522];
@(posedge clk);
#1;data_in = testData5[9523];
@(posedge clk);
#1;data_in = testData5[9524];
@(posedge clk);
#1;data_in = testData5[9525];
@(posedge clk);
#1;data_in = testData5[9526];
@(posedge clk);
#1;data_in = testData5[9527];
@(posedge clk);
#1;data_in = testData5[9528];
@(posedge clk);
#1;data_in = testData5[9529];
@(posedge clk);
#1;data_in = testData5[9530];
@(posedge clk);
#1;data_in = testData5[9531];
@(posedge clk);
#1;data_in = testData5[9532];
@(posedge clk);
#1;data_in = testData5[9533];
@(posedge clk);
#1;data_in = testData5[9534];
@(posedge clk);
#1;data_in = testData5[9535];
@(posedge clk);
#1;data_in = testData5[9536];
@(posedge clk);
#1;data_in = testData5[9537];
@(posedge clk);
#1;data_in = testData5[9538];
@(posedge clk);
#1;data_in = testData5[9539];
@(posedge clk);
#1;data_in = testData5[9540];
@(posedge clk);
#1;data_in = testData5[9541];
@(posedge clk);
#1;data_in = testData5[9542];
@(posedge clk);
#1;data_in = testData5[9543];
@(posedge clk);
#1;data_in = testData5[9544];
@(posedge clk);
#1;data_in = testData5[9545];
@(posedge clk);
#1;data_in = testData5[9546];
@(posedge clk);
#1;data_in = testData5[9547];
@(posedge clk);
#1;data_in = testData5[9548];
@(posedge clk);
#1;data_in = testData5[9549];
@(posedge clk);
#1;data_in = testData5[9550];
@(posedge clk);
#1;data_in = testData5[9551];
@(posedge clk);
#1;data_in = testData5[9552];
@(posedge clk);
#1;data_in = testData5[9553];
@(posedge clk);
#1;data_in = testData5[9554];
@(posedge clk);
#1;data_in = testData5[9555];
@(posedge clk);
#1;data_in = testData5[9556];
@(posedge clk);
#1;data_in = testData5[9557];
@(posedge clk);
#1;data_in = testData5[9558];
@(posedge clk);
#1;data_in = testData5[9559];
@(posedge clk);
#1;data_in = testData5[9560];
@(posedge clk);
#1;data_in = testData5[9561];
@(posedge clk);
#1;data_in = testData5[9562];
@(posedge clk);
#1;data_in = testData5[9563];
@(posedge clk);
#1;data_in = testData5[9564];
@(posedge clk);
#1;data_in = testData5[9565];
@(posedge clk);
#1;data_in = testData5[9566];
@(posedge clk);
#1;data_in = testData5[9567];
@(posedge clk);
#1;data_in = testData5[9568];
@(posedge clk);
#1;data_in = testData5[9569];
@(posedge clk);
#1;data_in = testData5[9570];
@(posedge clk);
#1;data_in = testData5[9571];
@(posedge clk);
#1;data_in = testData5[9572];
@(posedge clk);
#1;data_in = testData5[9573];
@(posedge clk);
#1;data_in = testData5[9574];
@(posedge clk);
#1;data_in = testData5[9575];
@(posedge clk);
#1;data_in = testData5[9576];
@(posedge clk);
#1;data_in = testData5[9577];
@(posedge clk);
#1;data_in = testData5[9578];
@(posedge clk);
#1;data_in = testData5[9579];
@(posedge clk);
#1;data_in = testData5[9580];
@(posedge clk);
#1;data_in = testData5[9581];
@(posedge clk);
#1;data_in = testData5[9582];
@(posedge clk);
#1;data_in = testData5[9583];
@(posedge clk);
#1;data_in = testData5[9584];
@(posedge clk);
#1;data_in = testData5[9585];
@(posedge clk);
#1;data_in = testData5[9586];
@(posedge clk);
#1;data_in = testData5[9587];
@(posedge clk);
#1;data_in = testData5[9588];
@(posedge clk);
#1;data_in = testData5[9589];
@(posedge clk);
#1;data_in = testData5[9590];
@(posedge clk);
#1;data_in = testData5[9591];
@(posedge clk);
#1;data_in = testData5[9592];
@(posedge clk);
#1;data_in = testData5[9593];
@(posedge clk);
#1;data_in = testData5[9594];
@(posedge clk);
#1;data_in = testData5[9595];
@(posedge clk);
#1;data_in = testData5[9596];
@(posedge clk);
#1;data_in = testData5[9597];
@(posedge clk);
#1;data_in = testData5[9598];
@(posedge clk);
#1;data_in = testData5[9599];
@(posedge clk);
#1;data_in = testData5[9600];
@(posedge clk);
#1;data_in = testData5[9601];
@(posedge clk);
#1;data_in = testData5[9602];
@(posedge clk);
#1;data_in = testData5[9603];
@(posedge clk);
#1;data_in = testData5[9604];
@(posedge clk);
#1;data_in = testData5[9605];
@(posedge clk);
#1;data_in = testData5[9606];
@(posedge clk);
#1;data_in = testData5[9607];
@(posedge clk);
#1;data_in = testData5[9608];
@(posedge clk);
#1;data_in = testData5[9609];
@(posedge clk);
#1;data_in = testData5[9610];
@(posedge clk);
#1;data_in = testData5[9611];
@(posedge clk);
#1;data_in = testData5[9612];
@(posedge clk);
#1;data_in = testData5[9613];
@(posedge clk);
#1;data_in = testData5[9614];
@(posedge clk);
#1;data_in = testData5[9615];
@(posedge clk);
#1;data_in = testData5[9616];
@(posedge clk);
#1;data_in = testData5[9617];
@(posedge clk);
#1;data_in = testData5[9618];
@(posedge clk);
#1;data_in = testData5[9619];
@(posedge clk);
#1;data_in = testData5[9620];
@(posedge clk);
#1;data_in = testData5[9621];
@(posedge clk);
#1;data_in = testData5[9622];
@(posedge clk);
#1;data_in = testData5[9623];
@(posedge clk);
#1;data_in = testData5[9624];
@(posedge clk);
#1;data_in = testData5[9625];
@(posedge clk);
#1;data_in = testData5[9626];
@(posedge clk);
#1;data_in = testData5[9627];
@(posedge clk);
#1;data_in = testData5[9628];
@(posedge clk);
#1;data_in = testData5[9629];
@(posedge clk);
#1;data_in = testData5[9630];
@(posedge clk);
#1;data_in = testData5[9631];
@(posedge clk);
#1;data_in = testData5[9632];
@(posedge clk);
#1;data_in = testData5[9633];
@(posedge clk);
#1;data_in = testData5[9634];
@(posedge clk);
#1;data_in = testData5[9635];
@(posedge clk);
#1;data_in = testData5[9636];
@(posedge clk);
#1;data_in = testData5[9637];
@(posedge clk);
#1;data_in = testData5[9638];
@(posedge clk);
#1;data_in = testData5[9639];
@(posedge clk);
#1;data_in = testData5[9640];
@(posedge clk);
#1;data_in = testData5[9641];
@(posedge clk);
#1;data_in = testData5[9642];
@(posedge clk);
#1;data_in = testData5[9643];
@(posedge clk);
#1;data_in = testData5[9644];
@(posedge clk);
#1;data_in = testData5[9645];
@(posedge clk);
#1;data_in = testData5[9646];
@(posedge clk);
#1;data_in = testData5[9647];
@(posedge clk);
#1;data_in = testData5[9648];
@(posedge clk);
#1;data_in = testData5[9649];
@(posedge clk);
#1;data_in = testData5[9650];
@(posedge clk);
#1;data_in = testData5[9651];
@(posedge clk);
#1;data_in = testData5[9652];
@(posedge clk);
#1;data_in = testData5[9653];
@(posedge clk);
#1;data_in = testData5[9654];
@(posedge clk);
#1;data_in = testData5[9655];
@(posedge clk);
#1;data_in = testData5[9656];
@(posedge clk);
#1;data_in = testData5[9657];
@(posedge clk);
#1;data_in = testData5[9658];
@(posedge clk);
#1;data_in = testData5[9659];
@(posedge clk);
#1;data_in = testData5[9660];
@(posedge clk);
#1;data_in = testData5[9661];
@(posedge clk);
#1;data_in = testData5[9662];
@(posedge clk);
#1;data_in = testData5[9663];
@(posedge clk);
#1;data_in = testData5[9664];
@(posedge clk);
#1;data_in = testData5[9665];
@(posedge clk);
#1;data_in = testData5[9666];
@(posedge clk);
#1;data_in = testData5[9667];
@(posedge clk);
#1;data_in = testData5[9668];
@(posedge clk);
#1;data_in = testData5[9669];
@(posedge clk);
#1;data_in = testData5[9670];
@(posedge clk);
#1;data_in = testData5[9671];
@(posedge clk);
#1;data_in = testData5[9672];
@(posedge clk);
#1;data_in = testData5[9673];
@(posedge clk);
#1;data_in = testData5[9674];
@(posedge clk);
#1;data_in = testData5[9675];
@(posedge clk);
#1;data_in = testData5[9676];
@(posedge clk);
#1;data_in = testData5[9677];
@(posedge clk);
#1;data_in = testData5[9678];
@(posedge clk);
#1;data_in = testData5[9679];
@(posedge clk);
#1;data_in = testData5[9680];
@(posedge clk);
#1;data_in = testData5[9681];
@(posedge clk);
#1;data_in = testData5[9682];
@(posedge clk);
#1;data_in = testData5[9683];
@(posedge clk);
#1;data_in = testData5[9684];
@(posedge clk);
#1;data_in = testData5[9685];
@(posedge clk);
#1;data_in = testData5[9686];
@(posedge clk);
#1;data_in = testData5[9687];
@(posedge clk);
#1;data_in = testData5[9688];
@(posedge clk);
#1;data_in = testData5[9689];
@(posedge clk);
#1;data_in = testData5[9690];
@(posedge clk);
#1;data_in = testData5[9691];
@(posedge clk);
#1;data_in = testData5[9692];
@(posedge clk);
#1;data_in = testData5[9693];
@(posedge clk);
#1;data_in = testData5[9694];
@(posedge clk);
#1;data_in = testData5[9695];
@(posedge clk);
#1;data_in = testData5[9696];
@(posedge clk);
#1;data_in = testData5[9697];
@(posedge clk);
#1;data_in = testData5[9698];
@(posedge clk);
#1;data_in = testData5[9699];
@(posedge clk);
#1;data_in = testData5[9700];
@(posedge clk);
#1;data_in = testData5[9701];
@(posedge clk);
#1;data_in = testData5[9702];
@(posedge clk);
#1;data_in = testData5[9703];
@(posedge clk);
#1;data_in = testData5[9704];
@(posedge clk);
#1;data_in = testData5[9705];
@(posedge clk);
#1;data_in = testData5[9706];
@(posedge clk);
#1;data_in = testData5[9707];
@(posedge clk);
#1;data_in = testData5[9708];
@(posedge clk);
#1;data_in = testData5[9709];
@(posedge clk);
#1;data_in = testData5[9710];
@(posedge clk);
#1;data_in = testData5[9711];
@(posedge clk);
#1;data_in = testData5[9712];
@(posedge clk);
#1;data_in = testData5[9713];
@(posedge clk);
#1;data_in = testData5[9714];
@(posedge clk);
#1;data_in = testData5[9715];
@(posedge clk);
#1;data_in = testData5[9716];
@(posedge clk);
#1;data_in = testData5[9717];
@(posedge clk);
#1;data_in = testData5[9718];
@(posedge clk);
#1;data_in = testData5[9719];
@(posedge clk);
#1;data_in = testData5[9720];
@(posedge clk);
#1;data_in = testData5[9721];
@(posedge clk);
#1;data_in = testData5[9722];
@(posedge clk);
#1;data_in = testData5[9723];
@(posedge clk);
#1;data_in = testData5[9724];
@(posedge clk);
#1;data_in = testData5[9725];
@(posedge clk);
#1;data_in = testData5[9726];
@(posedge clk);
#1;data_in = testData5[9727];
@(posedge clk);
#1;data_in = testData5[9728];
@(posedge clk);
#1;data_in = testData5[9729];
@(posedge clk);
#1;data_in = testData5[9730];
@(posedge clk);
#1;data_in = testData5[9731];
@(posedge clk);
#1;data_in = testData5[9732];
@(posedge clk);
#1;data_in = testData5[9733];
@(posedge clk);
#1;data_in = testData5[9734];
@(posedge clk);
#1;data_in = testData5[9735];
@(posedge clk);
#1;data_in = testData5[9736];
@(posedge clk);
#1;data_in = testData5[9737];
@(posedge clk);
#1;data_in = testData5[9738];
@(posedge clk);
#1;data_in = testData5[9739];
@(posedge clk);
#1;data_in = testData5[9740];
@(posedge clk);
#1;data_in = testData5[9741];
@(posedge clk);
#1;data_in = testData5[9742];
@(posedge clk);
#1;data_in = testData5[9743];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[9744]; 
@(posedge clk);
#1;data_in = testData5[9745];
@(posedge clk);
#1;data_in = testData5[9746];
@(posedge clk);
#1;data_in = testData5[9747];
@(posedge clk);
#1;data_in = testData5[9748];
@(posedge clk);
#1;data_in = testData5[9749];
@(posedge clk);
#1;data_in = testData5[9750];
@(posedge clk);
#1;data_in = testData5[9751];
@(posedge clk);
#1;data_in = testData5[9752];
@(posedge clk);
#1;data_in = testData5[9753];
@(posedge clk);
#1;data_in = testData5[9754];
@(posedge clk);
#1;data_in = testData5[9755];
@(posedge clk);
#1;data_in = testData5[9756];
@(posedge clk);
#1;data_in = testData5[9757];
@(posedge clk);
#1;data_in = testData5[9758];
@(posedge clk);
#1;data_in = testData5[9759];
@(posedge clk);
#1;data_in = testData5[9760];
@(posedge clk);
#1;data_in = testData5[9761];
@(posedge clk);
#1;data_in = testData5[9762];
@(posedge clk);
#1;data_in = testData5[9763];
@(posedge clk);
#1;data_in = testData5[9764];
@(posedge clk);
#1;data_in = testData5[9765];
@(posedge clk);
#1;data_in = testData5[9766];
@(posedge clk);
#1;data_in = testData5[9767];
@(posedge clk);
#1;data_in = testData5[9768];
@(posedge clk);
#1;data_in = testData5[9769];
@(posedge clk);
#1;data_in = testData5[9770];
@(posedge clk);
#1;data_in = testData5[9771];
@(posedge clk);
#1;data_in = testData5[9772];
@(posedge clk);
#1;data_in = testData5[9773];
@(posedge clk);
#1;data_in = testData5[9774];
@(posedge clk);
#1;data_in = testData5[9775];
@(posedge clk);
#1;data_in = testData5[9776];
@(posedge clk);
#1;data_in = testData5[9777];
@(posedge clk);
#1;data_in = testData5[9778];
@(posedge clk);
#1;data_in = testData5[9779];
@(posedge clk);
#1;data_in = testData5[9780];
@(posedge clk);
#1;data_in = testData5[9781];
@(posedge clk);
#1;data_in = testData5[9782];
@(posedge clk);
#1;data_in = testData5[9783];
@(posedge clk);
#1;data_in = testData5[9784];
@(posedge clk);
#1;data_in = testData5[9785];
@(posedge clk);
#1;data_in = testData5[9786];
@(posedge clk);
#1;data_in = testData5[9787];
@(posedge clk);
#1;data_in = testData5[9788];
@(posedge clk);
#1;data_in = testData5[9789];
@(posedge clk);
#1;data_in = testData5[9790];
@(posedge clk);
#1;data_in = testData5[9791];
@(posedge clk);
#1;data_in = testData5[9792];
@(posedge clk);
#1;data_in = testData5[9793];
@(posedge clk);
#1;data_in = testData5[9794];
@(posedge clk);
#1;data_in = testData5[9795];
@(posedge clk);
#1;data_in = testData5[9796];
@(posedge clk);
#1;data_in = testData5[9797];
@(posedge clk);
#1;data_in = testData5[9798];
@(posedge clk);
#1;data_in = testData5[9799];
@(posedge clk);
#1;data_in = testData5[9800];
@(posedge clk);
#1;data_in = testData5[9801];
@(posedge clk);
#1;data_in = testData5[9802];
@(posedge clk);
#1;data_in = testData5[9803];
@(posedge clk);
#1;data_in = testData5[9804];
@(posedge clk);
#1;data_in = testData5[9805];
@(posedge clk);
#1;data_in = testData5[9806];
@(posedge clk);
#1;data_in = testData5[9807];
@(posedge clk);
#1;data_in = testData5[9808];
@(posedge clk);
#1;data_in = testData5[9809];
@(posedge clk);
#1;data_in = testData5[9810];
@(posedge clk);
#1;data_in = testData5[9811];
@(posedge clk);
#1;data_in = testData5[9812];
@(posedge clk);
#1;data_in = testData5[9813];
@(posedge clk);
#1;data_in = testData5[9814];
@(posedge clk);
#1;data_in = testData5[9815];
@(posedge clk);
#1;data_in = testData5[9816];
@(posedge clk);
#1;data_in = testData5[9817];
@(posedge clk);
#1;data_in = testData5[9818];
@(posedge clk);
#1;data_in = testData5[9819];
@(posedge clk);
#1;data_in = testData5[9820];
@(posedge clk);
#1;data_in = testData5[9821];
@(posedge clk);
#1;data_in = testData5[9822];
@(posedge clk);
#1;data_in = testData5[9823];
@(posedge clk);
#1;data_in = testData5[9824];
@(posedge clk);
#1;data_in = testData5[9825];
@(posedge clk);
#1;data_in = testData5[9826];
@(posedge clk);
#1;data_in = testData5[9827];
@(posedge clk);
#1;data_in = testData5[9828];
@(posedge clk);
#1;data_in = testData5[9829];
@(posedge clk);
#1;data_in = testData5[9830];
@(posedge clk);
#1;data_in = testData5[9831];
@(posedge clk);
#1;data_in = testData5[9832];
@(posedge clk);
#1;data_in = testData5[9833];
@(posedge clk);
#1;data_in = testData5[9834];
@(posedge clk);
#1;data_in = testData5[9835];
@(posedge clk);
#1;data_in = testData5[9836];
@(posedge clk);
#1;data_in = testData5[9837];
@(posedge clk);
#1;data_in = testData5[9838];
@(posedge clk);
#1;data_in = testData5[9839];
@(posedge clk);
#1;data_in = testData5[9840];
@(posedge clk);
#1;data_in = testData5[9841];
@(posedge clk);
#1;data_in = testData5[9842];
@(posedge clk);
#1;data_in = testData5[9843];
@(posedge clk);
#1;data_in = testData5[9844];
@(posedge clk);
#1;data_in = testData5[9845];
@(posedge clk);
#1;data_in = testData5[9846];
@(posedge clk);
#1;data_in = testData5[9847];
@(posedge clk);
#1;data_in = testData5[9848];
@(posedge clk);
#1;data_in = testData5[9849];
@(posedge clk);
#1;data_in = testData5[9850];
@(posedge clk);
#1;data_in = testData5[9851];
@(posedge clk);
#1;data_in = testData5[9852];
@(posedge clk);
#1;data_in = testData5[9853];
@(posedge clk);
#1;data_in = testData5[9854];
@(posedge clk);
#1;data_in = testData5[9855];
@(posedge clk);
#1;data_in = testData5[9856];
@(posedge clk);
#1;data_in = testData5[9857];
@(posedge clk);
#1;data_in = testData5[9858];
@(posedge clk);
#1;data_in = testData5[9859];
@(posedge clk);
#1;data_in = testData5[9860];
@(posedge clk);
#1;data_in = testData5[9861];
@(posedge clk);
#1;data_in = testData5[9862];
@(posedge clk);
#1;data_in = testData5[9863];
@(posedge clk);
#1;data_in = testData5[9864];
@(posedge clk);
#1;data_in = testData5[9865];
@(posedge clk);
#1;data_in = testData5[9866];
@(posedge clk);
#1;data_in = testData5[9867];
@(posedge clk);
#1;data_in = testData5[9868];
@(posedge clk);
#1;data_in = testData5[9869];
@(posedge clk);
#1;data_in = testData5[9870];
@(posedge clk);
#1;data_in = testData5[9871];
@(posedge clk);
#1;data_in = testData5[9872];
@(posedge clk);
#1;data_in = testData5[9873];
@(posedge clk);
#1;data_in = testData5[9874];
@(posedge clk);
#1;data_in = testData5[9875];
@(posedge clk);
#1;data_in = testData5[9876];
@(posedge clk);
#1;data_in = testData5[9877];
@(posedge clk);
#1;data_in = testData5[9878];
@(posedge clk);
#1;data_in = testData5[9879];
@(posedge clk);
#1;data_in = testData5[9880];
@(posedge clk);
#1;data_in = testData5[9881];
@(posedge clk);
#1;data_in = testData5[9882];
@(posedge clk);
#1;data_in = testData5[9883];
@(posedge clk);
#1;data_in = testData5[9884];
@(posedge clk);
#1;data_in = testData5[9885];
@(posedge clk);
#1;data_in = testData5[9886];
@(posedge clk);
#1;data_in = testData5[9887];
@(posedge clk);
#1;data_in = testData5[9888];
@(posedge clk);
#1;data_in = testData5[9889];
@(posedge clk);
#1;data_in = testData5[9890];
@(posedge clk);
#1;data_in = testData5[9891];
@(posedge clk);
#1;data_in = testData5[9892];
@(posedge clk);
#1;data_in = testData5[9893];
@(posedge clk);
#1;data_in = testData5[9894];
@(posedge clk);
#1;data_in = testData5[9895];
@(posedge clk);
#1;data_in = testData5[9896];
@(posedge clk);
#1;data_in = testData5[9897];
@(posedge clk);
#1;data_in = testData5[9898];
@(posedge clk);
#1;data_in = testData5[9899];
@(posedge clk);
#1;data_in = testData5[9900];
@(posedge clk);
#1;data_in = testData5[9901];
@(posedge clk);
#1;data_in = testData5[9902];
@(posedge clk);
#1;data_in = testData5[9903];
@(posedge clk);
#1;data_in = testData5[9904];
@(posedge clk);
#1;data_in = testData5[9905];
@(posedge clk);
#1;data_in = testData5[9906];
@(posedge clk);
#1;data_in = testData5[9907];
@(posedge clk);
#1;data_in = testData5[9908];
@(posedge clk);
#1;data_in = testData5[9909];
@(posedge clk);
#1;data_in = testData5[9910];
@(posedge clk);
#1;data_in = testData5[9911];
@(posedge clk);
#1;data_in = testData5[9912];
@(posedge clk);
#1;data_in = testData5[9913];
@(posedge clk);
#1;data_in = testData5[9914];
@(posedge clk);
#1;data_in = testData5[9915];
@(posedge clk);
#1;data_in = testData5[9916];
@(posedge clk);
#1;data_in = testData5[9917];
@(posedge clk);
#1;data_in = testData5[9918];
@(posedge clk);
#1;data_in = testData5[9919];
@(posedge clk);
#1;data_in = testData5[9920];
@(posedge clk);
#1;data_in = testData5[9921];
@(posedge clk);
#1;data_in = testData5[9922];
@(posedge clk);
#1;data_in = testData5[9923];
@(posedge clk);
#1;data_in = testData5[9924];
@(posedge clk);
#1;data_in = testData5[9925];
@(posedge clk);
#1;data_in = testData5[9926];
@(posedge clk);
#1;data_in = testData5[9927];
@(posedge clk);
#1;data_in = testData5[9928];
@(posedge clk);
#1;data_in = testData5[9929];
@(posedge clk);
#1;data_in = testData5[9930];
@(posedge clk);
#1;data_in = testData5[9931];
@(posedge clk);
#1;data_in = testData5[9932];
@(posedge clk);
#1;data_in = testData5[9933];
@(posedge clk);
#1;data_in = testData5[9934];
@(posedge clk);
#1;data_in = testData5[9935];
@(posedge clk);
#1;data_in = testData5[9936];
@(posedge clk);
#1;data_in = testData5[9937];
@(posedge clk);
#1;data_in = testData5[9938];
@(posedge clk);
#1;data_in = testData5[9939];
@(posedge clk);
#1;data_in = testData5[9940];
@(posedge clk);
#1;data_in = testData5[9941];
@(posedge clk);
#1;data_in = testData5[9942];
@(posedge clk);
#1;data_in = testData5[9943];
@(posedge clk);
#1;data_in = testData5[9944];
@(posedge clk);
#1;data_in = testData5[9945];
@(posedge clk);
#1;data_in = testData5[9946];
@(posedge clk);
#1;data_in = testData5[9947];
@(posedge clk);
#1;data_in = testData5[9948];
@(posedge clk);
#1;data_in = testData5[9949];
@(posedge clk);
#1;data_in = testData5[9950];
@(posedge clk);
#1;data_in = testData5[9951];
@(posedge clk);
#1;data_in = testData5[9952];
@(posedge clk);
#1;data_in = testData5[9953];
@(posedge clk);
#1;data_in = testData5[9954];
@(posedge clk);
#1;data_in = testData5[9955];
@(posedge clk);
#1;data_in = testData5[9956];
@(posedge clk);
#1;data_in = testData5[9957];
@(posedge clk);
#1;data_in = testData5[9958];
@(posedge clk);
#1;data_in = testData5[9959];
@(posedge clk);
#1;data_in = testData5[9960];
@(posedge clk);
#1;data_in = testData5[9961];
@(posedge clk);
#1;data_in = testData5[9962];
@(posedge clk);
#1;data_in = testData5[9963];
@(posedge clk);
#1;data_in = testData5[9964];
@(posedge clk);
#1;data_in = testData5[9965];
@(posedge clk);
#1;data_in = testData5[9966];
@(posedge clk);
#1;data_in = testData5[9967];
@(posedge clk);
#1;data_in = testData5[9968];
@(posedge clk);
#1;data_in = testData5[9969];
@(posedge clk);
#1;data_in = testData5[9970];
@(posedge clk);
#1;data_in = testData5[9971];
@(posedge clk);
#1;data_in = testData5[9972];
@(posedge clk);
#1;data_in = testData5[9973];
@(posedge clk);
#1;data_in = testData5[9974];
@(posedge clk);
#1;data_in = testData5[9975];
@(posedge clk);
#1;data_in = testData5[9976];
@(posedge clk);
#1;data_in = testData5[9977];
@(posedge clk);
#1;data_in = testData5[9978];
@(posedge clk);
#1;data_in = testData5[9979];
@(posedge clk);
#1;data_in = testData5[9980];
@(posedge clk);
#1;data_in = testData5[9981];
@(posedge clk);
#1;data_in = testData5[9982];
@(posedge clk);
#1;data_in = testData5[9983];
@(posedge clk);
#1;data_in = testData5[9984];
@(posedge clk);
#1;data_in = testData5[9985];
@(posedge clk);
#1;data_in = testData5[9986];
@(posedge clk);
#1;data_in = testData5[9987];
@(posedge clk);
#1;data_in = testData5[9988];
@(posedge clk);
#1;data_in = testData5[9989];
@(posedge clk);
#1;data_in = testData5[9990];
@(posedge clk);
#1;data_in = testData5[9991];
@(posedge clk);
#1;data_in = testData5[9992];
@(posedge clk);
#1;data_in = testData5[9993];
@(posedge clk);
#1;data_in = testData5[9994];
@(posedge clk);
#1;data_in = testData5[9995];
@(posedge clk);
#1;data_in = testData5[9996];
@(posedge clk);
#1;data_in = testData5[9997];
@(posedge clk);
#1;data_in = testData5[9998];
@(posedge clk);
#1;data_in = testData5[9999];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[10000]; 
@(posedge clk);
#1;data_in = testData5[10001];
@(posedge clk);
#1;data_in = testData5[10002];
@(posedge clk);
#1;data_in = testData5[10003];
@(posedge clk);
#1;data_in = testData5[10004];
@(posedge clk);
#1;data_in = testData5[10005];
@(posedge clk);
#1;data_in = testData5[10006];
@(posedge clk);
#1;data_in = testData5[10007];
@(posedge clk);
#1;data_in = testData5[10008];
@(posedge clk);
#1;data_in = testData5[10009];
@(posedge clk);
#1;data_in = testData5[10010];
@(posedge clk);
#1;data_in = testData5[10011];
@(posedge clk);
#1;data_in = testData5[10012];
@(posedge clk);
#1;data_in = testData5[10013];
@(posedge clk);
#1;data_in = testData5[10014];
@(posedge clk);
#1;data_in = testData5[10015];
@(posedge clk);
#1;data_in = testData5[10016];
@(posedge clk);
#1;data_in = testData5[10017];
@(posedge clk);
#1;data_in = testData5[10018];
@(posedge clk);
#1;data_in = testData5[10019];
@(posedge clk);
#1;data_in = testData5[10020];
@(posedge clk);
#1;data_in = testData5[10021];
@(posedge clk);
#1;data_in = testData5[10022];
@(posedge clk);
#1;data_in = testData5[10023];
@(posedge clk);
#1;data_in = testData5[10024];
@(posedge clk);
#1;data_in = testData5[10025];
@(posedge clk);
#1;data_in = testData5[10026];
@(posedge clk);
#1;data_in = testData5[10027];
@(posedge clk);
#1;data_in = testData5[10028];
@(posedge clk);
#1;data_in = testData5[10029];
@(posedge clk);
#1;data_in = testData5[10030];
@(posedge clk);
#1;data_in = testData5[10031];
@(posedge clk);
#1;data_in = testData5[10032];
@(posedge clk);
#1;data_in = testData5[10033];
@(posedge clk);
#1;data_in = testData5[10034];
@(posedge clk);
#1;data_in = testData5[10035];
@(posedge clk);
#1;data_in = testData5[10036];
@(posedge clk);
#1;data_in = testData5[10037];
@(posedge clk);
#1;data_in = testData5[10038];
@(posedge clk);
#1;data_in = testData5[10039];
@(posedge clk);
#1;data_in = testData5[10040];
@(posedge clk);
#1;data_in = testData5[10041];
@(posedge clk);
#1;data_in = testData5[10042];
@(posedge clk);
#1;data_in = testData5[10043];
@(posedge clk);
#1;data_in = testData5[10044];
@(posedge clk);
#1;data_in = testData5[10045];
@(posedge clk);
#1;data_in = testData5[10046];
@(posedge clk);
#1;data_in = testData5[10047];
@(posedge clk);
#1;data_in = testData5[10048];
@(posedge clk);
#1;data_in = testData5[10049];
@(posedge clk);
#1;data_in = testData5[10050];
@(posedge clk);
#1;data_in = testData5[10051];
@(posedge clk);
#1;data_in = testData5[10052];
@(posedge clk);
#1;data_in = testData5[10053];
@(posedge clk);
#1;data_in = testData5[10054];
@(posedge clk);
#1;data_in = testData5[10055];
@(posedge clk);
#1;data_in = testData5[10056];
@(posedge clk);
#1;data_in = testData5[10057];
@(posedge clk);
#1;data_in = testData5[10058];
@(posedge clk);
#1;data_in = testData5[10059];
@(posedge clk);
#1;data_in = testData5[10060];
@(posedge clk);
#1;data_in = testData5[10061];
@(posedge clk);
#1;data_in = testData5[10062];
@(posedge clk);
#1;data_in = testData5[10063];
@(posedge clk);
#1;data_in = testData5[10064];
@(posedge clk);
#1;data_in = testData5[10065];
@(posedge clk);
#1;data_in = testData5[10066];
@(posedge clk);
#1;data_in = testData5[10067];
@(posedge clk);
#1;data_in = testData5[10068];
@(posedge clk);
#1;data_in = testData5[10069];
@(posedge clk);
#1;data_in = testData5[10070];
@(posedge clk);
#1;data_in = testData5[10071];
@(posedge clk);
#1;data_in = testData5[10072];
@(posedge clk);
#1;data_in = testData5[10073];
@(posedge clk);
#1;data_in = testData5[10074];
@(posedge clk);
#1;data_in = testData5[10075];
@(posedge clk);
#1;data_in = testData5[10076];
@(posedge clk);
#1;data_in = testData5[10077];
@(posedge clk);
#1;data_in = testData5[10078];
@(posedge clk);
#1;data_in = testData5[10079];
@(posedge clk);
#1;data_in = testData5[10080];
@(posedge clk);
#1;data_in = testData5[10081];
@(posedge clk);
#1;data_in = testData5[10082];
@(posedge clk);
#1;data_in = testData5[10083];
@(posedge clk);
#1;data_in = testData5[10084];
@(posedge clk);
#1;data_in = testData5[10085];
@(posedge clk);
#1;data_in = testData5[10086];
@(posedge clk);
#1;data_in = testData5[10087];
@(posedge clk);
#1;data_in = testData5[10088];
@(posedge clk);
#1;data_in = testData5[10089];
@(posedge clk);
#1;data_in = testData5[10090];
@(posedge clk);
#1;data_in = testData5[10091];
@(posedge clk);
#1;data_in = testData5[10092];
@(posedge clk);
#1;data_in = testData5[10093];
@(posedge clk);
#1;data_in = testData5[10094];
@(posedge clk);
#1;data_in = testData5[10095];
@(posedge clk);
#1;data_in = testData5[10096];
@(posedge clk);
#1;data_in = testData5[10097];
@(posedge clk);
#1;data_in = testData5[10098];
@(posedge clk);
#1;data_in = testData5[10099];
@(posedge clk);
#1;data_in = testData5[10100];
@(posedge clk);
#1;data_in = testData5[10101];
@(posedge clk);
#1;data_in = testData5[10102];
@(posedge clk);
#1;data_in = testData5[10103];
@(posedge clk);
#1;data_in = testData5[10104];
@(posedge clk);
#1;data_in = testData5[10105];
@(posedge clk);
#1;data_in = testData5[10106];
@(posedge clk);
#1;data_in = testData5[10107];
@(posedge clk);
#1;data_in = testData5[10108];
@(posedge clk);
#1;data_in = testData5[10109];
@(posedge clk);
#1;data_in = testData5[10110];
@(posedge clk);
#1;data_in = testData5[10111];
@(posedge clk);
#1;data_in = testData5[10112];
@(posedge clk);
#1;data_in = testData5[10113];
@(posedge clk);
#1;data_in = testData5[10114];
@(posedge clk);
#1;data_in = testData5[10115];
@(posedge clk);
#1;data_in = testData5[10116];
@(posedge clk);
#1;data_in = testData5[10117];
@(posedge clk);
#1;data_in = testData5[10118];
@(posedge clk);
#1;data_in = testData5[10119];
@(posedge clk);
#1;data_in = testData5[10120];
@(posedge clk);
#1;data_in = testData5[10121];
@(posedge clk);
#1;data_in = testData5[10122];
@(posedge clk);
#1;data_in = testData5[10123];
@(posedge clk);
#1;data_in = testData5[10124];
@(posedge clk);
#1;data_in = testData5[10125];
@(posedge clk);
#1;data_in = testData5[10126];
@(posedge clk);
#1;data_in = testData5[10127];
@(posedge clk);
#1;data_in = testData5[10128];
@(posedge clk);
#1;data_in = testData5[10129];
@(posedge clk);
#1;data_in = testData5[10130];
@(posedge clk);
#1;data_in = testData5[10131];
@(posedge clk);
#1;data_in = testData5[10132];
@(posedge clk);
#1;data_in = testData5[10133];
@(posedge clk);
#1;data_in = testData5[10134];
@(posedge clk);
#1;data_in = testData5[10135];
@(posedge clk);
#1;data_in = testData5[10136];
@(posedge clk);
#1;data_in = testData5[10137];
@(posedge clk);
#1;data_in = testData5[10138];
@(posedge clk);
#1;data_in = testData5[10139];
@(posedge clk);
#1;data_in = testData5[10140];
@(posedge clk);
#1;data_in = testData5[10141];
@(posedge clk);
#1;data_in = testData5[10142];
@(posedge clk);
#1;data_in = testData5[10143];
@(posedge clk);
#1;data_in = testData5[10144];
@(posedge clk);
#1;data_in = testData5[10145];
@(posedge clk);
#1;data_in = testData5[10146];
@(posedge clk);
#1;data_in = testData5[10147];
@(posedge clk);
#1;data_in = testData5[10148];
@(posedge clk);
#1;data_in = testData5[10149];
@(posedge clk);
#1;data_in = testData5[10150];
@(posedge clk);
#1;data_in = testData5[10151];
@(posedge clk);
#1;data_in = testData5[10152];
@(posedge clk);
#1;data_in = testData5[10153];
@(posedge clk);
#1;data_in = testData5[10154];
@(posedge clk);
#1;data_in = testData5[10155];
@(posedge clk);
#1;data_in = testData5[10156];
@(posedge clk);
#1;data_in = testData5[10157];
@(posedge clk);
#1;data_in = testData5[10158];
@(posedge clk);
#1;data_in = testData5[10159];
@(posedge clk);
#1;data_in = testData5[10160];
@(posedge clk);
#1;data_in = testData5[10161];
@(posedge clk);
#1;data_in = testData5[10162];
@(posedge clk);
#1;data_in = testData5[10163];
@(posedge clk);
#1;data_in = testData5[10164];
@(posedge clk);
#1;data_in = testData5[10165];
@(posedge clk);
#1;data_in = testData5[10166];
@(posedge clk);
#1;data_in = testData5[10167];
@(posedge clk);
#1;data_in = testData5[10168];
@(posedge clk);
#1;data_in = testData5[10169];
@(posedge clk);
#1;data_in = testData5[10170];
@(posedge clk);
#1;data_in = testData5[10171];
@(posedge clk);
#1;data_in = testData5[10172];
@(posedge clk);
#1;data_in = testData5[10173];
@(posedge clk);
#1;data_in = testData5[10174];
@(posedge clk);
#1;data_in = testData5[10175];
@(posedge clk);
#1;data_in = testData5[10176];
@(posedge clk);
#1;data_in = testData5[10177];
@(posedge clk);
#1;data_in = testData5[10178];
@(posedge clk);
#1;data_in = testData5[10179];
@(posedge clk);
#1;data_in = testData5[10180];
@(posedge clk);
#1;data_in = testData5[10181];
@(posedge clk);
#1;data_in = testData5[10182];
@(posedge clk);
#1;data_in = testData5[10183];
@(posedge clk);
#1;data_in = testData5[10184];
@(posedge clk);
#1;data_in = testData5[10185];
@(posedge clk);
#1;data_in = testData5[10186];
@(posedge clk);
#1;data_in = testData5[10187];
@(posedge clk);
#1;data_in = testData5[10188];
@(posedge clk);
#1;data_in = testData5[10189];
@(posedge clk);
#1;data_in = testData5[10190];
@(posedge clk);
#1;data_in = testData5[10191];
@(posedge clk);
#1;data_in = testData5[10192];
@(posedge clk);
#1;data_in = testData5[10193];
@(posedge clk);
#1;data_in = testData5[10194];
@(posedge clk);
#1;data_in = testData5[10195];
@(posedge clk);
#1;data_in = testData5[10196];
@(posedge clk);
#1;data_in = testData5[10197];
@(posedge clk);
#1;data_in = testData5[10198];
@(posedge clk);
#1;data_in = testData5[10199];
@(posedge clk);
#1;data_in = testData5[10200];
@(posedge clk);
#1;data_in = testData5[10201];
@(posedge clk);
#1;data_in = testData5[10202];
@(posedge clk);
#1;data_in = testData5[10203];
@(posedge clk);
#1;data_in = testData5[10204];
@(posedge clk);
#1;data_in = testData5[10205];
@(posedge clk);
#1;data_in = testData5[10206];
@(posedge clk);
#1;data_in = testData5[10207];
@(posedge clk);
#1;data_in = testData5[10208];
@(posedge clk);
#1;data_in = testData5[10209];
@(posedge clk);
#1;data_in = testData5[10210];
@(posedge clk);
#1;data_in = testData5[10211];
@(posedge clk);
#1;data_in = testData5[10212];
@(posedge clk);
#1;data_in = testData5[10213];
@(posedge clk);
#1;data_in = testData5[10214];
@(posedge clk);
#1;data_in = testData5[10215];
@(posedge clk);
#1;data_in = testData5[10216];
@(posedge clk);
#1;data_in = testData5[10217];
@(posedge clk);
#1;data_in = testData5[10218];
@(posedge clk);
#1;data_in = testData5[10219];
@(posedge clk);
#1;data_in = testData5[10220];
@(posedge clk);
#1;data_in = testData5[10221];
@(posedge clk);
#1;data_in = testData5[10222];
@(posedge clk);
#1;data_in = testData5[10223];
@(posedge clk);
#1;data_in = testData5[10224];
@(posedge clk);
#1;data_in = testData5[10225];
@(posedge clk);
#1;data_in = testData5[10226];
@(posedge clk);
#1;data_in = testData5[10227];
@(posedge clk);
#1;data_in = testData5[10228];
@(posedge clk);
#1;data_in = testData5[10229];
@(posedge clk);
#1;data_in = testData5[10230];
@(posedge clk);
#1;data_in = testData5[10231];
@(posedge clk);
#1;data_in = testData5[10232];
@(posedge clk);
#1;data_in = testData5[10233];
@(posedge clk);
#1;data_in = testData5[10234];
@(posedge clk);
#1;data_in = testData5[10235];
@(posedge clk);
#1;data_in = testData5[10236];
@(posedge clk);
#1;data_in = testData5[10237];
@(posedge clk);
#1;data_in = testData5[10238];
@(posedge clk);
#1;data_in = testData5[10239];
@(posedge clk);
#1;data_in = testData5[10240];
@(posedge clk);
#1;data_in = testData5[10241];
@(posedge clk);
#1;data_in = testData5[10242];
@(posedge clk);
#1;data_in = testData5[10243];
@(posedge clk);
#1;data_in = testData5[10244];
@(posedge clk);
#1;data_in = testData5[10245];
@(posedge clk);
#1;data_in = testData5[10246];
@(posedge clk);
#1;data_in = testData5[10247];
@(posedge clk);
#1;data_in = testData5[10248];
@(posedge clk);
#1;data_in = testData5[10249];
@(posedge clk);
#1;data_in = testData5[10250];
@(posedge clk);
#1;data_in = testData5[10251];
@(posedge clk);
#1;data_in = testData5[10252];
@(posedge clk);
#1;data_in = testData5[10253];
@(posedge clk);
#1;data_in = testData5[10254];
@(posedge clk);
#1;data_in = testData5[10255];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[10256]; 
@(posedge clk);
#1;data_in = testData5[10257];
@(posedge clk);
#1;data_in = testData5[10258];
@(posedge clk);
#1;data_in = testData5[10259];
@(posedge clk);
#1;data_in = testData5[10260];
@(posedge clk);
#1;data_in = testData5[10261];
@(posedge clk);
#1;data_in = testData5[10262];
@(posedge clk);
#1;data_in = testData5[10263];
@(posedge clk);
#1;data_in = testData5[10264];
@(posedge clk);
#1;data_in = testData5[10265];
@(posedge clk);
#1;data_in = testData5[10266];
@(posedge clk);
#1;data_in = testData5[10267];
@(posedge clk);
#1;data_in = testData5[10268];
@(posedge clk);
#1;data_in = testData5[10269];
@(posedge clk);
#1;data_in = testData5[10270];
@(posedge clk);
#1;data_in = testData5[10271];
@(posedge clk);
#1;data_in = testData5[10272];
@(posedge clk);
#1;data_in = testData5[10273];
@(posedge clk);
#1;data_in = testData5[10274];
@(posedge clk);
#1;data_in = testData5[10275];
@(posedge clk);
#1;data_in = testData5[10276];
@(posedge clk);
#1;data_in = testData5[10277];
@(posedge clk);
#1;data_in = testData5[10278];
@(posedge clk);
#1;data_in = testData5[10279];
@(posedge clk);
#1;data_in = testData5[10280];
@(posedge clk);
#1;data_in = testData5[10281];
@(posedge clk);
#1;data_in = testData5[10282];
@(posedge clk);
#1;data_in = testData5[10283];
@(posedge clk);
#1;data_in = testData5[10284];
@(posedge clk);
#1;data_in = testData5[10285];
@(posedge clk);
#1;data_in = testData5[10286];
@(posedge clk);
#1;data_in = testData5[10287];
@(posedge clk);
#1;data_in = testData5[10288];
@(posedge clk);
#1;data_in = testData5[10289];
@(posedge clk);
#1;data_in = testData5[10290];
@(posedge clk);
#1;data_in = testData5[10291];
@(posedge clk);
#1;data_in = testData5[10292];
@(posedge clk);
#1;data_in = testData5[10293];
@(posedge clk);
#1;data_in = testData5[10294];
@(posedge clk);
#1;data_in = testData5[10295];
@(posedge clk);
#1;data_in = testData5[10296];
@(posedge clk);
#1;data_in = testData5[10297];
@(posedge clk);
#1;data_in = testData5[10298];
@(posedge clk);
#1;data_in = testData5[10299];
@(posedge clk);
#1;data_in = testData5[10300];
@(posedge clk);
#1;data_in = testData5[10301];
@(posedge clk);
#1;data_in = testData5[10302];
@(posedge clk);
#1;data_in = testData5[10303];
@(posedge clk);
#1;data_in = testData5[10304];
@(posedge clk);
#1;data_in = testData5[10305];
@(posedge clk);
#1;data_in = testData5[10306];
@(posedge clk);
#1;data_in = testData5[10307];
@(posedge clk);
#1;data_in = testData5[10308];
@(posedge clk);
#1;data_in = testData5[10309];
@(posedge clk);
#1;data_in = testData5[10310];
@(posedge clk);
#1;data_in = testData5[10311];
@(posedge clk);
#1;data_in = testData5[10312];
@(posedge clk);
#1;data_in = testData5[10313];
@(posedge clk);
#1;data_in = testData5[10314];
@(posedge clk);
#1;data_in = testData5[10315];
@(posedge clk);
#1;data_in = testData5[10316];
@(posedge clk);
#1;data_in = testData5[10317];
@(posedge clk);
#1;data_in = testData5[10318];
@(posedge clk);
#1;data_in = testData5[10319];
@(posedge clk);
#1;data_in = testData5[10320];
@(posedge clk);
#1;data_in = testData5[10321];
@(posedge clk);
#1;data_in = testData5[10322];
@(posedge clk);
#1;data_in = testData5[10323];
@(posedge clk);
#1;data_in = testData5[10324];
@(posedge clk);
#1;data_in = testData5[10325];
@(posedge clk);
#1;data_in = testData5[10326];
@(posedge clk);
#1;data_in = testData5[10327];
@(posedge clk);
#1;data_in = testData5[10328];
@(posedge clk);
#1;data_in = testData5[10329];
@(posedge clk);
#1;data_in = testData5[10330];
@(posedge clk);
#1;data_in = testData5[10331];
@(posedge clk);
#1;data_in = testData5[10332];
@(posedge clk);
#1;data_in = testData5[10333];
@(posedge clk);
#1;data_in = testData5[10334];
@(posedge clk);
#1;data_in = testData5[10335];
@(posedge clk);
#1;data_in = testData5[10336];
@(posedge clk);
#1;data_in = testData5[10337];
@(posedge clk);
#1;data_in = testData5[10338];
@(posedge clk);
#1;data_in = testData5[10339];
@(posedge clk);
#1;data_in = testData5[10340];
@(posedge clk);
#1;data_in = testData5[10341];
@(posedge clk);
#1;data_in = testData5[10342];
@(posedge clk);
#1;data_in = testData5[10343];
@(posedge clk);
#1;data_in = testData5[10344];
@(posedge clk);
#1;data_in = testData5[10345];
@(posedge clk);
#1;data_in = testData5[10346];
@(posedge clk);
#1;data_in = testData5[10347];
@(posedge clk);
#1;data_in = testData5[10348];
@(posedge clk);
#1;data_in = testData5[10349];
@(posedge clk);
#1;data_in = testData5[10350];
@(posedge clk);
#1;data_in = testData5[10351];
@(posedge clk);
#1;data_in = testData5[10352];
@(posedge clk);
#1;data_in = testData5[10353];
@(posedge clk);
#1;data_in = testData5[10354];
@(posedge clk);
#1;data_in = testData5[10355];
@(posedge clk);
#1;data_in = testData5[10356];
@(posedge clk);
#1;data_in = testData5[10357];
@(posedge clk);
#1;data_in = testData5[10358];
@(posedge clk);
#1;data_in = testData5[10359];
@(posedge clk);
#1;data_in = testData5[10360];
@(posedge clk);
#1;data_in = testData5[10361];
@(posedge clk);
#1;data_in = testData5[10362];
@(posedge clk);
#1;data_in = testData5[10363];
@(posedge clk);
#1;data_in = testData5[10364];
@(posedge clk);
#1;data_in = testData5[10365];
@(posedge clk);
#1;data_in = testData5[10366];
@(posedge clk);
#1;data_in = testData5[10367];
@(posedge clk);
#1;data_in = testData5[10368];
@(posedge clk);
#1;data_in = testData5[10369];
@(posedge clk);
#1;data_in = testData5[10370];
@(posedge clk);
#1;data_in = testData5[10371];
@(posedge clk);
#1;data_in = testData5[10372];
@(posedge clk);
#1;data_in = testData5[10373];
@(posedge clk);
#1;data_in = testData5[10374];
@(posedge clk);
#1;data_in = testData5[10375];
@(posedge clk);
#1;data_in = testData5[10376];
@(posedge clk);
#1;data_in = testData5[10377];
@(posedge clk);
#1;data_in = testData5[10378];
@(posedge clk);
#1;data_in = testData5[10379];
@(posedge clk);
#1;data_in = testData5[10380];
@(posedge clk);
#1;data_in = testData5[10381];
@(posedge clk);
#1;data_in = testData5[10382];
@(posedge clk);
#1;data_in = testData5[10383];
@(posedge clk);
#1;data_in = testData5[10384];
@(posedge clk);
#1;data_in = testData5[10385];
@(posedge clk);
#1;data_in = testData5[10386];
@(posedge clk);
#1;data_in = testData5[10387];
@(posedge clk);
#1;data_in = testData5[10388];
@(posedge clk);
#1;data_in = testData5[10389];
@(posedge clk);
#1;data_in = testData5[10390];
@(posedge clk);
#1;data_in = testData5[10391];
@(posedge clk);
#1;data_in = testData5[10392];
@(posedge clk);
#1;data_in = testData5[10393];
@(posedge clk);
#1;data_in = testData5[10394];
@(posedge clk);
#1;data_in = testData5[10395];
@(posedge clk);
#1;data_in = testData5[10396];
@(posedge clk);
#1;data_in = testData5[10397];
@(posedge clk);
#1;data_in = testData5[10398];
@(posedge clk);
#1;data_in = testData5[10399];
@(posedge clk);
#1;data_in = testData5[10400];
@(posedge clk);
#1;data_in = testData5[10401];
@(posedge clk);
#1;data_in = testData5[10402];
@(posedge clk);
#1;data_in = testData5[10403];
@(posedge clk);
#1;data_in = testData5[10404];
@(posedge clk);
#1;data_in = testData5[10405];
@(posedge clk);
#1;data_in = testData5[10406];
@(posedge clk);
#1;data_in = testData5[10407];
@(posedge clk);
#1;data_in = testData5[10408];
@(posedge clk);
#1;data_in = testData5[10409];
@(posedge clk);
#1;data_in = testData5[10410];
@(posedge clk);
#1;data_in = testData5[10411];
@(posedge clk);
#1;data_in = testData5[10412];
@(posedge clk);
#1;data_in = testData5[10413];
@(posedge clk);
#1;data_in = testData5[10414];
@(posedge clk);
#1;data_in = testData5[10415];
@(posedge clk);
#1;data_in = testData5[10416];
@(posedge clk);
#1;data_in = testData5[10417];
@(posedge clk);
#1;data_in = testData5[10418];
@(posedge clk);
#1;data_in = testData5[10419];
@(posedge clk);
#1;data_in = testData5[10420];
@(posedge clk);
#1;data_in = testData5[10421];
@(posedge clk);
#1;data_in = testData5[10422];
@(posedge clk);
#1;data_in = testData5[10423];
@(posedge clk);
#1;data_in = testData5[10424];
@(posedge clk);
#1;data_in = testData5[10425];
@(posedge clk);
#1;data_in = testData5[10426];
@(posedge clk);
#1;data_in = testData5[10427];
@(posedge clk);
#1;data_in = testData5[10428];
@(posedge clk);
#1;data_in = testData5[10429];
@(posedge clk);
#1;data_in = testData5[10430];
@(posedge clk);
#1;data_in = testData5[10431];
@(posedge clk);
#1;data_in = testData5[10432];
@(posedge clk);
#1;data_in = testData5[10433];
@(posedge clk);
#1;data_in = testData5[10434];
@(posedge clk);
#1;data_in = testData5[10435];
@(posedge clk);
#1;data_in = testData5[10436];
@(posedge clk);
#1;data_in = testData5[10437];
@(posedge clk);
#1;data_in = testData5[10438];
@(posedge clk);
#1;data_in = testData5[10439];
@(posedge clk);
#1;data_in = testData5[10440];
@(posedge clk);
#1;data_in = testData5[10441];
@(posedge clk);
#1;data_in = testData5[10442];
@(posedge clk);
#1;data_in = testData5[10443];
@(posedge clk);
#1;data_in = testData5[10444];
@(posedge clk);
#1;data_in = testData5[10445];
@(posedge clk);
#1;data_in = testData5[10446];
@(posedge clk);
#1;data_in = testData5[10447];
@(posedge clk);
#1;data_in = testData5[10448];
@(posedge clk);
#1;data_in = testData5[10449];
@(posedge clk);
#1;data_in = testData5[10450];
@(posedge clk);
#1;data_in = testData5[10451];
@(posedge clk);
#1;data_in = testData5[10452];
@(posedge clk);
#1;data_in = testData5[10453];
@(posedge clk);
#1;data_in = testData5[10454];
@(posedge clk);
#1;data_in = testData5[10455];
@(posedge clk);
#1;data_in = testData5[10456];
@(posedge clk);
#1;data_in = testData5[10457];
@(posedge clk);
#1;data_in = testData5[10458];
@(posedge clk);
#1;data_in = testData5[10459];
@(posedge clk);
#1;data_in = testData5[10460];
@(posedge clk);
#1;data_in = testData5[10461];
@(posedge clk);
#1;data_in = testData5[10462];
@(posedge clk);
#1;data_in = testData5[10463];
@(posedge clk);
#1;data_in = testData5[10464];
@(posedge clk);
#1;data_in = testData5[10465];
@(posedge clk);
#1;data_in = testData5[10466];
@(posedge clk);
#1;data_in = testData5[10467];
@(posedge clk);
#1;data_in = testData5[10468];
@(posedge clk);
#1;data_in = testData5[10469];
@(posedge clk);
#1;data_in = testData5[10470];
@(posedge clk);
#1;data_in = testData5[10471];
@(posedge clk);
#1;data_in = testData5[10472];
@(posedge clk);
#1;data_in = testData5[10473];
@(posedge clk);
#1;data_in = testData5[10474];
@(posedge clk);
#1;data_in = testData5[10475];
@(posedge clk);
#1;data_in = testData5[10476];
@(posedge clk);
#1;data_in = testData5[10477];
@(posedge clk);
#1;data_in = testData5[10478];
@(posedge clk);
#1;data_in = testData5[10479];
@(posedge clk);
#1;data_in = testData5[10480];
@(posedge clk);
#1;data_in = testData5[10481];
@(posedge clk);
#1;data_in = testData5[10482];
@(posedge clk);
#1;data_in = testData5[10483];
@(posedge clk);
#1;data_in = testData5[10484];
@(posedge clk);
#1;data_in = testData5[10485];
@(posedge clk);
#1;data_in = testData5[10486];
@(posedge clk);
#1;data_in = testData5[10487];
@(posedge clk);
#1;data_in = testData5[10488];
@(posedge clk);
#1;data_in = testData5[10489];
@(posedge clk);
#1;data_in = testData5[10490];
@(posedge clk);
#1;data_in = testData5[10491];
@(posedge clk);
#1;data_in = testData5[10492];
@(posedge clk);
#1;data_in = testData5[10493];
@(posedge clk);
#1;data_in = testData5[10494];
@(posedge clk);
#1;data_in = testData5[10495];
@(posedge clk);
#1;data_in = testData5[10496];
@(posedge clk);
#1;data_in = testData5[10497];
@(posedge clk);
#1;data_in = testData5[10498];
@(posedge clk);
#1;data_in = testData5[10499];
@(posedge clk);
#1;data_in = testData5[10500];
@(posedge clk);
#1;data_in = testData5[10501];
@(posedge clk);
#1;data_in = testData5[10502];
@(posedge clk);
#1;data_in = testData5[10503];
@(posedge clk);
#1;data_in = testData5[10504];
@(posedge clk);
#1;data_in = testData5[10505];
@(posedge clk);
#1;data_in = testData5[10506];
@(posedge clk);
#1;data_in = testData5[10507];
@(posedge clk);
#1;data_in = testData5[10508];
@(posedge clk);
#1;data_in = testData5[10509];
@(posedge clk);
#1;data_in = testData5[10510];
@(posedge clk);
#1;data_in = testData5[10511];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[10512]; 
@(posedge clk);
#1;data_in = testData5[10513];
@(posedge clk);
#1;data_in = testData5[10514];
@(posedge clk);
#1;data_in = testData5[10515];
@(posedge clk);
#1;data_in = testData5[10516];
@(posedge clk);
#1;data_in = testData5[10517];
@(posedge clk);
#1;data_in = testData5[10518];
@(posedge clk);
#1;data_in = testData5[10519];
@(posedge clk);
#1;data_in = testData5[10520];
@(posedge clk);
#1;data_in = testData5[10521];
@(posedge clk);
#1;data_in = testData5[10522];
@(posedge clk);
#1;data_in = testData5[10523];
@(posedge clk);
#1;data_in = testData5[10524];
@(posedge clk);
#1;data_in = testData5[10525];
@(posedge clk);
#1;data_in = testData5[10526];
@(posedge clk);
#1;data_in = testData5[10527];
@(posedge clk);
#1;data_in = testData5[10528];
@(posedge clk);
#1;data_in = testData5[10529];
@(posedge clk);
#1;data_in = testData5[10530];
@(posedge clk);
#1;data_in = testData5[10531];
@(posedge clk);
#1;data_in = testData5[10532];
@(posedge clk);
#1;data_in = testData5[10533];
@(posedge clk);
#1;data_in = testData5[10534];
@(posedge clk);
#1;data_in = testData5[10535];
@(posedge clk);
#1;data_in = testData5[10536];
@(posedge clk);
#1;data_in = testData5[10537];
@(posedge clk);
#1;data_in = testData5[10538];
@(posedge clk);
#1;data_in = testData5[10539];
@(posedge clk);
#1;data_in = testData5[10540];
@(posedge clk);
#1;data_in = testData5[10541];
@(posedge clk);
#1;data_in = testData5[10542];
@(posedge clk);
#1;data_in = testData5[10543];
@(posedge clk);
#1;data_in = testData5[10544];
@(posedge clk);
#1;data_in = testData5[10545];
@(posedge clk);
#1;data_in = testData5[10546];
@(posedge clk);
#1;data_in = testData5[10547];
@(posedge clk);
#1;data_in = testData5[10548];
@(posedge clk);
#1;data_in = testData5[10549];
@(posedge clk);
#1;data_in = testData5[10550];
@(posedge clk);
#1;data_in = testData5[10551];
@(posedge clk);
#1;data_in = testData5[10552];
@(posedge clk);
#1;data_in = testData5[10553];
@(posedge clk);
#1;data_in = testData5[10554];
@(posedge clk);
#1;data_in = testData5[10555];
@(posedge clk);
#1;data_in = testData5[10556];
@(posedge clk);
#1;data_in = testData5[10557];
@(posedge clk);
#1;data_in = testData5[10558];
@(posedge clk);
#1;data_in = testData5[10559];
@(posedge clk);
#1;data_in = testData5[10560];
@(posedge clk);
#1;data_in = testData5[10561];
@(posedge clk);
#1;data_in = testData5[10562];
@(posedge clk);
#1;data_in = testData5[10563];
@(posedge clk);
#1;data_in = testData5[10564];
@(posedge clk);
#1;data_in = testData5[10565];
@(posedge clk);
#1;data_in = testData5[10566];
@(posedge clk);
#1;data_in = testData5[10567];
@(posedge clk);
#1;data_in = testData5[10568];
@(posedge clk);
#1;data_in = testData5[10569];
@(posedge clk);
#1;data_in = testData5[10570];
@(posedge clk);
#1;data_in = testData5[10571];
@(posedge clk);
#1;data_in = testData5[10572];
@(posedge clk);
#1;data_in = testData5[10573];
@(posedge clk);
#1;data_in = testData5[10574];
@(posedge clk);
#1;data_in = testData5[10575];
@(posedge clk);
#1;data_in = testData5[10576];
@(posedge clk);
#1;data_in = testData5[10577];
@(posedge clk);
#1;data_in = testData5[10578];
@(posedge clk);
#1;data_in = testData5[10579];
@(posedge clk);
#1;data_in = testData5[10580];
@(posedge clk);
#1;data_in = testData5[10581];
@(posedge clk);
#1;data_in = testData5[10582];
@(posedge clk);
#1;data_in = testData5[10583];
@(posedge clk);
#1;data_in = testData5[10584];
@(posedge clk);
#1;data_in = testData5[10585];
@(posedge clk);
#1;data_in = testData5[10586];
@(posedge clk);
#1;data_in = testData5[10587];
@(posedge clk);
#1;data_in = testData5[10588];
@(posedge clk);
#1;data_in = testData5[10589];
@(posedge clk);
#1;data_in = testData5[10590];
@(posedge clk);
#1;data_in = testData5[10591];
@(posedge clk);
#1;data_in = testData5[10592];
@(posedge clk);
#1;data_in = testData5[10593];
@(posedge clk);
#1;data_in = testData5[10594];
@(posedge clk);
#1;data_in = testData5[10595];
@(posedge clk);
#1;data_in = testData5[10596];
@(posedge clk);
#1;data_in = testData5[10597];
@(posedge clk);
#1;data_in = testData5[10598];
@(posedge clk);
#1;data_in = testData5[10599];
@(posedge clk);
#1;data_in = testData5[10600];
@(posedge clk);
#1;data_in = testData5[10601];
@(posedge clk);
#1;data_in = testData5[10602];
@(posedge clk);
#1;data_in = testData5[10603];
@(posedge clk);
#1;data_in = testData5[10604];
@(posedge clk);
#1;data_in = testData5[10605];
@(posedge clk);
#1;data_in = testData5[10606];
@(posedge clk);
#1;data_in = testData5[10607];
@(posedge clk);
#1;data_in = testData5[10608];
@(posedge clk);
#1;data_in = testData5[10609];
@(posedge clk);
#1;data_in = testData5[10610];
@(posedge clk);
#1;data_in = testData5[10611];
@(posedge clk);
#1;data_in = testData5[10612];
@(posedge clk);
#1;data_in = testData5[10613];
@(posedge clk);
#1;data_in = testData5[10614];
@(posedge clk);
#1;data_in = testData5[10615];
@(posedge clk);
#1;data_in = testData5[10616];
@(posedge clk);
#1;data_in = testData5[10617];
@(posedge clk);
#1;data_in = testData5[10618];
@(posedge clk);
#1;data_in = testData5[10619];
@(posedge clk);
#1;data_in = testData5[10620];
@(posedge clk);
#1;data_in = testData5[10621];
@(posedge clk);
#1;data_in = testData5[10622];
@(posedge clk);
#1;data_in = testData5[10623];
@(posedge clk);
#1;data_in = testData5[10624];
@(posedge clk);
#1;data_in = testData5[10625];
@(posedge clk);
#1;data_in = testData5[10626];
@(posedge clk);
#1;data_in = testData5[10627];
@(posedge clk);
#1;data_in = testData5[10628];
@(posedge clk);
#1;data_in = testData5[10629];
@(posedge clk);
#1;data_in = testData5[10630];
@(posedge clk);
#1;data_in = testData5[10631];
@(posedge clk);
#1;data_in = testData5[10632];
@(posedge clk);
#1;data_in = testData5[10633];
@(posedge clk);
#1;data_in = testData5[10634];
@(posedge clk);
#1;data_in = testData5[10635];
@(posedge clk);
#1;data_in = testData5[10636];
@(posedge clk);
#1;data_in = testData5[10637];
@(posedge clk);
#1;data_in = testData5[10638];
@(posedge clk);
#1;data_in = testData5[10639];
@(posedge clk);
#1;data_in = testData5[10640];
@(posedge clk);
#1;data_in = testData5[10641];
@(posedge clk);
#1;data_in = testData5[10642];
@(posedge clk);
#1;data_in = testData5[10643];
@(posedge clk);
#1;data_in = testData5[10644];
@(posedge clk);
#1;data_in = testData5[10645];
@(posedge clk);
#1;data_in = testData5[10646];
@(posedge clk);
#1;data_in = testData5[10647];
@(posedge clk);
#1;data_in = testData5[10648];
@(posedge clk);
#1;data_in = testData5[10649];
@(posedge clk);
#1;data_in = testData5[10650];
@(posedge clk);
#1;data_in = testData5[10651];
@(posedge clk);
#1;data_in = testData5[10652];
@(posedge clk);
#1;data_in = testData5[10653];
@(posedge clk);
#1;data_in = testData5[10654];
@(posedge clk);
#1;data_in = testData5[10655];
@(posedge clk);
#1;data_in = testData5[10656];
@(posedge clk);
#1;data_in = testData5[10657];
@(posedge clk);
#1;data_in = testData5[10658];
@(posedge clk);
#1;data_in = testData5[10659];
@(posedge clk);
#1;data_in = testData5[10660];
@(posedge clk);
#1;data_in = testData5[10661];
@(posedge clk);
#1;data_in = testData5[10662];
@(posedge clk);
#1;data_in = testData5[10663];
@(posedge clk);
#1;data_in = testData5[10664];
@(posedge clk);
#1;data_in = testData5[10665];
@(posedge clk);
#1;data_in = testData5[10666];
@(posedge clk);
#1;data_in = testData5[10667];
@(posedge clk);
#1;data_in = testData5[10668];
@(posedge clk);
#1;data_in = testData5[10669];
@(posedge clk);
#1;data_in = testData5[10670];
@(posedge clk);
#1;data_in = testData5[10671];
@(posedge clk);
#1;data_in = testData5[10672];
@(posedge clk);
#1;data_in = testData5[10673];
@(posedge clk);
#1;data_in = testData5[10674];
@(posedge clk);
#1;data_in = testData5[10675];
@(posedge clk);
#1;data_in = testData5[10676];
@(posedge clk);
#1;data_in = testData5[10677];
@(posedge clk);
#1;data_in = testData5[10678];
@(posedge clk);
#1;data_in = testData5[10679];
@(posedge clk);
#1;data_in = testData5[10680];
@(posedge clk);
#1;data_in = testData5[10681];
@(posedge clk);
#1;data_in = testData5[10682];
@(posedge clk);
#1;data_in = testData5[10683];
@(posedge clk);
#1;data_in = testData5[10684];
@(posedge clk);
#1;data_in = testData5[10685];
@(posedge clk);
#1;data_in = testData5[10686];
@(posedge clk);
#1;data_in = testData5[10687];
@(posedge clk);
#1;data_in = testData5[10688];
@(posedge clk);
#1;data_in = testData5[10689];
@(posedge clk);
#1;data_in = testData5[10690];
@(posedge clk);
#1;data_in = testData5[10691];
@(posedge clk);
#1;data_in = testData5[10692];
@(posedge clk);
#1;data_in = testData5[10693];
@(posedge clk);
#1;data_in = testData5[10694];
@(posedge clk);
#1;data_in = testData5[10695];
@(posedge clk);
#1;data_in = testData5[10696];
@(posedge clk);
#1;data_in = testData5[10697];
@(posedge clk);
#1;data_in = testData5[10698];
@(posedge clk);
#1;data_in = testData5[10699];
@(posedge clk);
#1;data_in = testData5[10700];
@(posedge clk);
#1;data_in = testData5[10701];
@(posedge clk);
#1;data_in = testData5[10702];
@(posedge clk);
#1;data_in = testData5[10703];
@(posedge clk);
#1;data_in = testData5[10704];
@(posedge clk);
#1;data_in = testData5[10705];
@(posedge clk);
#1;data_in = testData5[10706];
@(posedge clk);
#1;data_in = testData5[10707];
@(posedge clk);
#1;data_in = testData5[10708];
@(posedge clk);
#1;data_in = testData5[10709];
@(posedge clk);
#1;data_in = testData5[10710];
@(posedge clk);
#1;data_in = testData5[10711];
@(posedge clk);
#1;data_in = testData5[10712];
@(posedge clk);
#1;data_in = testData5[10713];
@(posedge clk);
#1;data_in = testData5[10714];
@(posedge clk);
#1;data_in = testData5[10715];
@(posedge clk);
#1;data_in = testData5[10716];
@(posedge clk);
#1;data_in = testData5[10717];
@(posedge clk);
#1;data_in = testData5[10718];
@(posedge clk);
#1;data_in = testData5[10719];
@(posedge clk);
#1;data_in = testData5[10720];
@(posedge clk);
#1;data_in = testData5[10721];
@(posedge clk);
#1;data_in = testData5[10722];
@(posedge clk);
#1;data_in = testData5[10723];
@(posedge clk);
#1;data_in = testData5[10724];
@(posedge clk);
#1;data_in = testData5[10725];
@(posedge clk);
#1;data_in = testData5[10726];
@(posedge clk);
#1;data_in = testData5[10727];
@(posedge clk);
#1;data_in = testData5[10728];
@(posedge clk);
#1;data_in = testData5[10729];
@(posedge clk);
#1;data_in = testData5[10730];
@(posedge clk);
#1;data_in = testData5[10731];
@(posedge clk);
#1;data_in = testData5[10732];
@(posedge clk);
#1;data_in = testData5[10733];
@(posedge clk);
#1;data_in = testData5[10734];
@(posedge clk);
#1;data_in = testData5[10735];
@(posedge clk);
#1;data_in = testData5[10736];
@(posedge clk);
#1;data_in = testData5[10737];
@(posedge clk);
#1;data_in = testData5[10738];
@(posedge clk);
#1;data_in = testData5[10739];
@(posedge clk);
#1;data_in = testData5[10740];
@(posedge clk);
#1;data_in = testData5[10741];
@(posedge clk);
#1;data_in = testData5[10742];
@(posedge clk);
#1;data_in = testData5[10743];
@(posedge clk);
#1;data_in = testData5[10744];
@(posedge clk);
#1;data_in = testData5[10745];
@(posedge clk);
#1;data_in = testData5[10746];
@(posedge clk);
#1;data_in = testData5[10747];
@(posedge clk);
#1;data_in = testData5[10748];
@(posedge clk);
#1;data_in = testData5[10749];
@(posedge clk);
#1;data_in = testData5[10750];
@(posedge clk);
#1;data_in = testData5[10751];
@(posedge clk);
#1;data_in = testData5[10752];
@(posedge clk);
#1;data_in = testData5[10753];
@(posedge clk);
#1;data_in = testData5[10754];
@(posedge clk);
#1;data_in = testData5[10755];
@(posedge clk);
#1;data_in = testData5[10756];
@(posedge clk);
#1;data_in = testData5[10757];
@(posedge clk);
#1;data_in = testData5[10758];
@(posedge clk);
#1;data_in = testData5[10759];
@(posedge clk);
#1;data_in = testData5[10760];
@(posedge clk);
#1;data_in = testData5[10761];
@(posedge clk);
#1;data_in = testData5[10762];
@(posedge clk);
#1;data_in = testData5[10763];
@(posedge clk);
#1;data_in = testData5[10764];
@(posedge clk);
#1;data_in = testData5[10765];
@(posedge clk);
#1;data_in = testData5[10766];
@(posedge clk);
#1;data_in = testData5[10767];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[10768]; 
@(posedge clk);
#1;data_in = testData5[10769];
@(posedge clk);
#1;data_in = testData5[10770];
@(posedge clk);
#1;data_in = testData5[10771];
@(posedge clk);
#1;data_in = testData5[10772];
@(posedge clk);
#1;data_in = testData5[10773];
@(posedge clk);
#1;data_in = testData5[10774];
@(posedge clk);
#1;data_in = testData5[10775];
@(posedge clk);
#1;data_in = testData5[10776];
@(posedge clk);
#1;data_in = testData5[10777];
@(posedge clk);
#1;data_in = testData5[10778];
@(posedge clk);
#1;data_in = testData5[10779];
@(posedge clk);
#1;data_in = testData5[10780];
@(posedge clk);
#1;data_in = testData5[10781];
@(posedge clk);
#1;data_in = testData5[10782];
@(posedge clk);
#1;data_in = testData5[10783];
@(posedge clk);
#1;data_in = testData5[10784];
@(posedge clk);
#1;data_in = testData5[10785];
@(posedge clk);
#1;data_in = testData5[10786];
@(posedge clk);
#1;data_in = testData5[10787];
@(posedge clk);
#1;data_in = testData5[10788];
@(posedge clk);
#1;data_in = testData5[10789];
@(posedge clk);
#1;data_in = testData5[10790];
@(posedge clk);
#1;data_in = testData5[10791];
@(posedge clk);
#1;data_in = testData5[10792];
@(posedge clk);
#1;data_in = testData5[10793];
@(posedge clk);
#1;data_in = testData5[10794];
@(posedge clk);
#1;data_in = testData5[10795];
@(posedge clk);
#1;data_in = testData5[10796];
@(posedge clk);
#1;data_in = testData5[10797];
@(posedge clk);
#1;data_in = testData5[10798];
@(posedge clk);
#1;data_in = testData5[10799];
@(posedge clk);
#1;data_in = testData5[10800];
@(posedge clk);
#1;data_in = testData5[10801];
@(posedge clk);
#1;data_in = testData5[10802];
@(posedge clk);
#1;data_in = testData5[10803];
@(posedge clk);
#1;data_in = testData5[10804];
@(posedge clk);
#1;data_in = testData5[10805];
@(posedge clk);
#1;data_in = testData5[10806];
@(posedge clk);
#1;data_in = testData5[10807];
@(posedge clk);
#1;data_in = testData5[10808];
@(posedge clk);
#1;data_in = testData5[10809];
@(posedge clk);
#1;data_in = testData5[10810];
@(posedge clk);
#1;data_in = testData5[10811];
@(posedge clk);
#1;data_in = testData5[10812];
@(posedge clk);
#1;data_in = testData5[10813];
@(posedge clk);
#1;data_in = testData5[10814];
@(posedge clk);
#1;data_in = testData5[10815];
@(posedge clk);
#1;data_in = testData5[10816];
@(posedge clk);
#1;data_in = testData5[10817];
@(posedge clk);
#1;data_in = testData5[10818];
@(posedge clk);
#1;data_in = testData5[10819];
@(posedge clk);
#1;data_in = testData5[10820];
@(posedge clk);
#1;data_in = testData5[10821];
@(posedge clk);
#1;data_in = testData5[10822];
@(posedge clk);
#1;data_in = testData5[10823];
@(posedge clk);
#1;data_in = testData5[10824];
@(posedge clk);
#1;data_in = testData5[10825];
@(posedge clk);
#1;data_in = testData5[10826];
@(posedge clk);
#1;data_in = testData5[10827];
@(posedge clk);
#1;data_in = testData5[10828];
@(posedge clk);
#1;data_in = testData5[10829];
@(posedge clk);
#1;data_in = testData5[10830];
@(posedge clk);
#1;data_in = testData5[10831];
@(posedge clk);
#1;data_in = testData5[10832];
@(posedge clk);
#1;data_in = testData5[10833];
@(posedge clk);
#1;data_in = testData5[10834];
@(posedge clk);
#1;data_in = testData5[10835];
@(posedge clk);
#1;data_in = testData5[10836];
@(posedge clk);
#1;data_in = testData5[10837];
@(posedge clk);
#1;data_in = testData5[10838];
@(posedge clk);
#1;data_in = testData5[10839];
@(posedge clk);
#1;data_in = testData5[10840];
@(posedge clk);
#1;data_in = testData5[10841];
@(posedge clk);
#1;data_in = testData5[10842];
@(posedge clk);
#1;data_in = testData5[10843];
@(posedge clk);
#1;data_in = testData5[10844];
@(posedge clk);
#1;data_in = testData5[10845];
@(posedge clk);
#1;data_in = testData5[10846];
@(posedge clk);
#1;data_in = testData5[10847];
@(posedge clk);
#1;data_in = testData5[10848];
@(posedge clk);
#1;data_in = testData5[10849];
@(posedge clk);
#1;data_in = testData5[10850];
@(posedge clk);
#1;data_in = testData5[10851];
@(posedge clk);
#1;data_in = testData5[10852];
@(posedge clk);
#1;data_in = testData5[10853];
@(posedge clk);
#1;data_in = testData5[10854];
@(posedge clk);
#1;data_in = testData5[10855];
@(posedge clk);
#1;data_in = testData5[10856];
@(posedge clk);
#1;data_in = testData5[10857];
@(posedge clk);
#1;data_in = testData5[10858];
@(posedge clk);
#1;data_in = testData5[10859];
@(posedge clk);
#1;data_in = testData5[10860];
@(posedge clk);
#1;data_in = testData5[10861];
@(posedge clk);
#1;data_in = testData5[10862];
@(posedge clk);
#1;data_in = testData5[10863];
@(posedge clk);
#1;data_in = testData5[10864];
@(posedge clk);
#1;data_in = testData5[10865];
@(posedge clk);
#1;data_in = testData5[10866];
@(posedge clk);
#1;data_in = testData5[10867];
@(posedge clk);
#1;data_in = testData5[10868];
@(posedge clk);
#1;data_in = testData5[10869];
@(posedge clk);
#1;data_in = testData5[10870];
@(posedge clk);
#1;data_in = testData5[10871];
@(posedge clk);
#1;data_in = testData5[10872];
@(posedge clk);
#1;data_in = testData5[10873];
@(posedge clk);
#1;data_in = testData5[10874];
@(posedge clk);
#1;data_in = testData5[10875];
@(posedge clk);
#1;data_in = testData5[10876];
@(posedge clk);
#1;data_in = testData5[10877];
@(posedge clk);
#1;data_in = testData5[10878];
@(posedge clk);
#1;data_in = testData5[10879];
@(posedge clk);
#1;data_in = testData5[10880];
@(posedge clk);
#1;data_in = testData5[10881];
@(posedge clk);
#1;data_in = testData5[10882];
@(posedge clk);
#1;data_in = testData5[10883];
@(posedge clk);
#1;data_in = testData5[10884];
@(posedge clk);
#1;data_in = testData5[10885];
@(posedge clk);
#1;data_in = testData5[10886];
@(posedge clk);
#1;data_in = testData5[10887];
@(posedge clk);
#1;data_in = testData5[10888];
@(posedge clk);
#1;data_in = testData5[10889];
@(posedge clk);
#1;data_in = testData5[10890];
@(posedge clk);
#1;data_in = testData5[10891];
@(posedge clk);
#1;data_in = testData5[10892];
@(posedge clk);
#1;data_in = testData5[10893];
@(posedge clk);
#1;data_in = testData5[10894];
@(posedge clk);
#1;data_in = testData5[10895];
@(posedge clk);
#1;data_in = testData5[10896];
@(posedge clk);
#1;data_in = testData5[10897];
@(posedge clk);
#1;data_in = testData5[10898];
@(posedge clk);
#1;data_in = testData5[10899];
@(posedge clk);
#1;data_in = testData5[10900];
@(posedge clk);
#1;data_in = testData5[10901];
@(posedge clk);
#1;data_in = testData5[10902];
@(posedge clk);
#1;data_in = testData5[10903];
@(posedge clk);
#1;data_in = testData5[10904];
@(posedge clk);
#1;data_in = testData5[10905];
@(posedge clk);
#1;data_in = testData5[10906];
@(posedge clk);
#1;data_in = testData5[10907];
@(posedge clk);
#1;data_in = testData5[10908];
@(posedge clk);
#1;data_in = testData5[10909];
@(posedge clk);
#1;data_in = testData5[10910];
@(posedge clk);
#1;data_in = testData5[10911];
@(posedge clk);
#1;data_in = testData5[10912];
@(posedge clk);
#1;data_in = testData5[10913];
@(posedge clk);
#1;data_in = testData5[10914];
@(posedge clk);
#1;data_in = testData5[10915];
@(posedge clk);
#1;data_in = testData5[10916];
@(posedge clk);
#1;data_in = testData5[10917];
@(posedge clk);
#1;data_in = testData5[10918];
@(posedge clk);
#1;data_in = testData5[10919];
@(posedge clk);
#1;data_in = testData5[10920];
@(posedge clk);
#1;data_in = testData5[10921];
@(posedge clk);
#1;data_in = testData5[10922];
@(posedge clk);
#1;data_in = testData5[10923];
@(posedge clk);
#1;data_in = testData5[10924];
@(posedge clk);
#1;data_in = testData5[10925];
@(posedge clk);
#1;data_in = testData5[10926];
@(posedge clk);
#1;data_in = testData5[10927];
@(posedge clk);
#1;data_in = testData5[10928];
@(posedge clk);
#1;data_in = testData5[10929];
@(posedge clk);
#1;data_in = testData5[10930];
@(posedge clk);
#1;data_in = testData5[10931];
@(posedge clk);
#1;data_in = testData5[10932];
@(posedge clk);
#1;data_in = testData5[10933];
@(posedge clk);
#1;data_in = testData5[10934];
@(posedge clk);
#1;data_in = testData5[10935];
@(posedge clk);
#1;data_in = testData5[10936];
@(posedge clk);
#1;data_in = testData5[10937];
@(posedge clk);
#1;data_in = testData5[10938];
@(posedge clk);
#1;data_in = testData5[10939];
@(posedge clk);
#1;data_in = testData5[10940];
@(posedge clk);
#1;data_in = testData5[10941];
@(posedge clk);
#1;data_in = testData5[10942];
@(posedge clk);
#1;data_in = testData5[10943];
@(posedge clk);
#1;data_in = testData5[10944];
@(posedge clk);
#1;data_in = testData5[10945];
@(posedge clk);
#1;data_in = testData5[10946];
@(posedge clk);
#1;data_in = testData5[10947];
@(posedge clk);
#1;data_in = testData5[10948];
@(posedge clk);
#1;data_in = testData5[10949];
@(posedge clk);
#1;data_in = testData5[10950];
@(posedge clk);
#1;data_in = testData5[10951];
@(posedge clk);
#1;data_in = testData5[10952];
@(posedge clk);
#1;data_in = testData5[10953];
@(posedge clk);
#1;data_in = testData5[10954];
@(posedge clk);
#1;data_in = testData5[10955];
@(posedge clk);
#1;data_in = testData5[10956];
@(posedge clk);
#1;data_in = testData5[10957];
@(posedge clk);
#1;data_in = testData5[10958];
@(posedge clk);
#1;data_in = testData5[10959];
@(posedge clk);
#1;data_in = testData5[10960];
@(posedge clk);
#1;data_in = testData5[10961];
@(posedge clk);
#1;data_in = testData5[10962];
@(posedge clk);
#1;data_in = testData5[10963];
@(posedge clk);
#1;data_in = testData5[10964];
@(posedge clk);
#1;data_in = testData5[10965];
@(posedge clk);
#1;data_in = testData5[10966];
@(posedge clk);
#1;data_in = testData5[10967];
@(posedge clk);
#1;data_in = testData5[10968];
@(posedge clk);
#1;data_in = testData5[10969];
@(posedge clk);
#1;data_in = testData5[10970];
@(posedge clk);
#1;data_in = testData5[10971];
@(posedge clk);
#1;data_in = testData5[10972];
@(posedge clk);
#1;data_in = testData5[10973];
@(posedge clk);
#1;data_in = testData5[10974];
@(posedge clk);
#1;data_in = testData5[10975];
@(posedge clk);
#1;data_in = testData5[10976];
@(posedge clk);
#1;data_in = testData5[10977];
@(posedge clk);
#1;data_in = testData5[10978];
@(posedge clk);
#1;data_in = testData5[10979];
@(posedge clk);
#1;data_in = testData5[10980];
@(posedge clk);
#1;data_in = testData5[10981];
@(posedge clk);
#1;data_in = testData5[10982];
@(posedge clk);
#1;data_in = testData5[10983];
@(posedge clk);
#1;data_in = testData5[10984];
@(posedge clk);
#1;data_in = testData5[10985];
@(posedge clk);
#1;data_in = testData5[10986];
@(posedge clk);
#1;data_in = testData5[10987];
@(posedge clk);
#1;data_in = testData5[10988];
@(posedge clk);
#1;data_in = testData5[10989];
@(posedge clk);
#1;data_in = testData5[10990];
@(posedge clk);
#1;data_in = testData5[10991];
@(posedge clk);
#1;data_in = testData5[10992];
@(posedge clk);
#1;data_in = testData5[10993];
@(posedge clk);
#1;data_in = testData5[10994];
@(posedge clk);
#1;data_in = testData5[10995];
@(posedge clk);
#1;data_in = testData5[10996];
@(posedge clk);
#1;data_in = testData5[10997];
@(posedge clk);
#1;data_in = testData5[10998];
@(posedge clk);
#1;data_in = testData5[10999];
@(posedge clk);
#1;data_in = testData5[11000];
@(posedge clk);
#1;data_in = testData5[11001];
@(posedge clk);
#1;data_in = testData5[11002];
@(posedge clk);
#1;data_in = testData5[11003];
@(posedge clk);
#1;data_in = testData5[11004];
@(posedge clk);
#1;data_in = testData5[11005];
@(posedge clk);
#1;data_in = testData5[11006];
@(posedge clk);
#1;data_in = testData5[11007];
@(posedge clk);
#1;data_in = testData5[11008];
@(posedge clk);
#1;data_in = testData5[11009];
@(posedge clk);
#1;data_in = testData5[11010];
@(posedge clk);
#1;data_in = testData5[11011];
@(posedge clk);
#1;data_in = testData5[11012];
@(posedge clk);
#1;data_in = testData5[11013];
@(posedge clk);
#1;data_in = testData5[11014];
@(posedge clk);
#1;data_in = testData5[11015];
@(posedge clk);
#1;data_in = testData5[11016];
@(posedge clk);
#1;data_in = testData5[11017];
@(posedge clk);
#1;data_in = testData5[11018];
@(posedge clk);
#1;data_in = testData5[11019];
@(posedge clk);
#1;data_in = testData5[11020];
@(posedge clk);
#1;data_in = testData5[11021];
@(posedge clk);
#1;data_in = testData5[11022];
@(posedge clk);
#1;data_in = testData5[11023];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[11024]; 
@(posedge clk);
#1;data_in = testData5[11025];
@(posedge clk);
#1;data_in = testData5[11026];
@(posedge clk);
#1;data_in = testData5[11027];
@(posedge clk);
#1;data_in = testData5[11028];
@(posedge clk);
#1;data_in = testData5[11029];
@(posedge clk);
#1;data_in = testData5[11030];
@(posedge clk);
#1;data_in = testData5[11031];
@(posedge clk);
#1;data_in = testData5[11032];
@(posedge clk);
#1;data_in = testData5[11033];
@(posedge clk);
#1;data_in = testData5[11034];
@(posedge clk);
#1;data_in = testData5[11035];
@(posedge clk);
#1;data_in = testData5[11036];
@(posedge clk);
#1;data_in = testData5[11037];
@(posedge clk);
#1;data_in = testData5[11038];
@(posedge clk);
#1;data_in = testData5[11039];
@(posedge clk);
#1;data_in = testData5[11040];
@(posedge clk);
#1;data_in = testData5[11041];
@(posedge clk);
#1;data_in = testData5[11042];
@(posedge clk);
#1;data_in = testData5[11043];
@(posedge clk);
#1;data_in = testData5[11044];
@(posedge clk);
#1;data_in = testData5[11045];
@(posedge clk);
#1;data_in = testData5[11046];
@(posedge clk);
#1;data_in = testData5[11047];
@(posedge clk);
#1;data_in = testData5[11048];
@(posedge clk);
#1;data_in = testData5[11049];
@(posedge clk);
#1;data_in = testData5[11050];
@(posedge clk);
#1;data_in = testData5[11051];
@(posedge clk);
#1;data_in = testData5[11052];
@(posedge clk);
#1;data_in = testData5[11053];
@(posedge clk);
#1;data_in = testData5[11054];
@(posedge clk);
#1;data_in = testData5[11055];
@(posedge clk);
#1;data_in = testData5[11056];
@(posedge clk);
#1;data_in = testData5[11057];
@(posedge clk);
#1;data_in = testData5[11058];
@(posedge clk);
#1;data_in = testData5[11059];
@(posedge clk);
#1;data_in = testData5[11060];
@(posedge clk);
#1;data_in = testData5[11061];
@(posedge clk);
#1;data_in = testData5[11062];
@(posedge clk);
#1;data_in = testData5[11063];
@(posedge clk);
#1;data_in = testData5[11064];
@(posedge clk);
#1;data_in = testData5[11065];
@(posedge clk);
#1;data_in = testData5[11066];
@(posedge clk);
#1;data_in = testData5[11067];
@(posedge clk);
#1;data_in = testData5[11068];
@(posedge clk);
#1;data_in = testData5[11069];
@(posedge clk);
#1;data_in = testData5[11070];
@(posedge clk);
#1;data_in = testData5[11071];
@(posedge clk);
#1;data_in = testData5[11072];
@(posedge clk);
#1;data_in = testData5[11073];
@(posedge clk);
#1;data_in = testData5[11074];
@(posedge clk);
#1;data_in = testData5[11075];
@(posedge clk);
#1;data_in = testData5[11076];
@(posedge clk);
#1;data_in = testData5[11077];
@(posedge clk);
#1;data_in = testData5[11078];
@(posedge clk);
#1;data_in = testData5[11079];
@(posedge clk);
#1;data_in = testData5[11080];
@(posedge clk);
#1;data_in = testData5[11081];
@(posedge clk);
#1;data_in = testData5[11082];
@(posedge clk);
#1;data_in = testData5[11083];
@(posedge clk);
#1;data_in = testData5[11084];
@(posedge clk);
#1;data_in = testData5[11085];
@(posedge clk);
#1;data_in = testData5[11086];
@(posedge clk);
#1;data_in = testData5[11087];
@(posedge clk);
#1;data_in = testData5[11088];
@(posedge clk);
#1;data_in = testData5[11089];
@(posedge clk);
#1;data_in = testData5[11090];
@(posedge clk);
#1;data_in = testData5[11091];
@(posedge clk);
#1;data_in = testData5[11092];
@(posedge clk);
#1;data_in = testData5[11093];
@(posedge clk);
#1;data_in = testData5[11094];
@(posedge clk);
#1;data_in = testData5[11095];
@(posedge clk);
#1;data_in = testData5[11096];
@(posedge clk);
#1;data_in = testData5[11097];
@(posedge clk);
#1;data_in = testData5[11098];
@(posedge clk);
#1;data_in = testData5[11099];
@(posedge clk);
#1;data_in = testData5[11100];
@(posedge clk);
#1;data_in = testData5[11101];
@(posedge clk);
#1;data_in = testData5[11102];
@(posedge clk);
#1;data_in = testData5[11103];
@(posedge clk);
#1;data_in = testData5[11104];
@(posedge clk);
#1;data_in = testData5[11105];
@(posedge clk);
#1;data_in = testData5[11106];
@(posedge clk);
#1;data_in = testData5[11107];
@(posedge clk);
#1;data_in = testData5[11108];
@(posedge clk);
#1;data_in = testData5[11109];
@(posedge clk);
#1;data_in = testData5[11110];
@(posedge clk);
#1;data_in = testData5[11111];
@(posedge clk);
#1;data_in = testData5[11112];
@(posedge clk);
#1;data_in = testData5[11113];
@(posedge clk);
#1;data_in = testData5[11114];
@(posedge clk);
#1;data_in = testData5[11115];
@(posedge clk);
#1;data_in = testData5[11116];
@(posedge clk);
#1;data_in = testData5[11117];
@(posedge clk);
#1;data_in = testData5[11118];
@(posedge clk);
#1;data_in = testData5[11119];
@(posedge clk);
#1;data_in = testData5[11120];
@(posedge clk);
#1;data_in = testData5[11121];
@(posedge clk);
#1;data_in = testData5[11122];
@(posedge clk);
#1;data_in = testData5[11123];
@(posedge clk);
#1;data_in = testData5[11124];
@(posedge clk);
#1;data_in = testData5[11125];
@(posedge clk);
#1;data_in = testData5[11126];
@(posedge clk);
#1;data_in = testData5[11127];
@(posedge clk);
#1;data_in = testData5[11128];
@(posedge clk);
#1;data_in = testData5[11129];
@(posedge clk);
#1;data_in = testData5[11130];
@(posedge clk);
#1;data_in = testData5[11131];
@(posedge clk);
#1;data_in = testData5[11132];
@(posedge clk);
#1;data_in = testData5[11133];
@(posedge clk);
#1;data_in = testData5[11134];
@(posedge clk);
#1;data_in = testData5[11135];
@(posedge clk);
#1;data_in = testData5[11136];
@(posedge clk);
#1;data_in = testData5[11137];
@(posedge clk);
#1;data_in = testData5[11138];
@(posedge clk);
#1;data_in = testData5[11139];
@(posedge clk);
#1;data_in = testData5[11140];
@(posedge clk);
#1;data_in = testData5[11141];
@(posedge clk);
#1;data_in = testData5[11142];
@(posedge clk);
#1;data_in = testData5[11143];
@(posedge clk);
#1;data_in = testData5[11144];
@(posedge clk);
#1;data_in = testData5[11145];
@(posedge clk);
#1;data_in = testData5[11146];
@(posedge clk);
#1;data_in = testData5[11147];
@(posedge clk);
#1;data_in = testData5[11148];
@(posedge clk);
#1;data_in = testData5[11149];
@(posedge clk);
#1;data_in = testData5[11150];
@(posedge clk);
#1;data_in = testData5[11151];
@(posedge clk);
#1;data_in = testData5[11152];
@(posedge clk);
#1;data_in = testData5[11153];
@(posedge clk);
#1;data_in = testData5[11154];
@(posedge clk);
#1;data_in = testData5[11155];
@(posedge clk);
#1;data_in = testData5[11156];
@(posedge clk);
#1;data_in = testData5[11157];
@(posedge clk);
#1;data_in = testData5[11158];
@(posedge clk);
#1;data_in = testData5[11159];
@(posedge clk);
#1;data_in = testData5[11160];
@(posedge clk);
#1;data_in = testData5[11161];
@(posedge clk);
#1;data_in = testData5[11162];
@(posedge clk);
#1;data_in = testData5[11163];
@(posedge clk);
#1;data_in = testData5[11164];
@(posedge clk);
#1;data_in = testData5[11165];
@(posedge clk);
#1;data_in = testData5[11166];
@(posedge clk);
#1;data_in = testData5[11167];
@(posedge clk);
#1;data_in = testData5[11168];
@(posedge clk);
#1;data_in = testData5[11169];
@(posedge clk);
#1;data_in = testData5[11170];
@(posedge clk);
#1;data_in = testData5[11171];
@(posedge clk);
#1;data_in = testData5[11172];
@(posedge clk);
#1;data_in = testData5[11173];
@(posedge clk);
#1;data_in = testData5[11174];
@(posedge clk);
#1;data_in = testData5[11175];
@(posedge clk);
#1;data_in = testData5[11176];
@(posedge clk);
#1;data_in = testData5[11177];
@(posedge clk);
#1;data_in = testData5[11178];
@(posedge clk);
#1;data_in = testData5[11179];
@(posedge clk);
#1;data_in = testData5[11180];
@(posedge clk);
#1;data_in = testData5[11181];
@(posedge clk);
#1;data_in = testData5[11182];
@(posedge clk);
#1;data_in = testData5[11183];
@(posedge clk);
#1;data_in = testData5[11184];
@(posedge clk);
#1;data_in = testData5[11185];
@(posedge clk);
#1;data_in = testData5[11186];
@(posedge clk);
#1;data_in = testData5[11187];
@(posedge clk);
#1;data_in = testData5[11188];
@(posedge clk);
#1;data_in = testData5[11189];
@(posedge clk);
#1;data_in = testData5[11190];
@(posedge clk);
#1;data_in = testData5[11191];
@(posedge clk);
#1;data_in = testData5[11192];
@(posedge clk);
#1;data_in = testData5[11193];
@(posedge clk);
#1;data_in = testData5[11194];
@(posedge clk);
#1;data_in = testData5[11195];
@(posedge clk);
#1;data_in = testData5[11196];
@(posedge clk);
#1;data_in = testData5[11197];
@(posedge clk);
#1;data_in = testData5[11198];
@(posedge clk);
#1;data_in = testData5[11199];
@(posedge clk);
#1;data_in = testData5[11200];
@(posedge clk);
#1;data_in = testData5[11201];
@(posedge clk);
#1;data_in = testData5[11202];
@(posedge clk);
#1;data_in = testData5[11203];
@(posedge clk);
#1;data_in = testData5[11204];
@(posedge clk);
#1;data_in = testData5[11205];
@(posedge clk);
#1;data_in = testData5[11206];
@(posedge clk);
#1;data_in = testData5[11207];
@(posedge clk);
#1;data_in = testData5[11208];
@(posedge clk);
#1;data_in = testData5[11209];
@(posedge clk);
#1;data_in = testData5[11210];
@(posedge clk);
#1;data_in = testData5[11211];
@(posedge clk);
#1;data_in = testData5[11212];
@(posedge clk);
#1;data_in = testData5[11213];
@(posedge clk);
#1;data_in = testData5[11214];
@(posedge clk);
#1;data_in = testData5[11215];
@(posedge clk);
#1;data_in = testData5[11216];
@(posedge clk);
#1;data_in = testData5[11217];
@(posedge clk);
#1;data_in = testData5[11218];
@(posedge clk);
#1;data_in = testData5[11219];
@(posedge clk);
#1;data_in = testData5[11220];
@(posedge clk);
#1;data_in = testData5[11221];
@(posedge clk);
#1;data_in = testData5[11222];
@(posedge clk);
#1;data_in = testData5[11223];
@(posedge clk);
#1;data_in = testData5[11224];
@(posedge clk);
#1;data_in = testData5[11225];
@(posedge clk);
#1;data_in = testData5[11226];
@(posedge clk);
#1;data_in = testData5[11227];
@(posedge clk);
#1;data_in = testData5[11228];
@(posedge clk);
#1;data_in = testData5[11229];
@(posedge clk);
#1;data_in = testData5[11230];
@(posedge clk);
#1;data_in = testData5[11231];
@(posedge clk);
#1;data_in = testData5[11232];
@(posedge clk);
#1;data_in = testData5[11233];
@(posedge clk);
#1;data_in = testData5[11234];
@(posedge clk);
#1;data_in = testData5[11235];
@(posedge clk);
#1;data_in = testData5[11236];
@(posedge clk);
#1;data_in = testData5[11237];
@(posedge clk);
#1;data_in = testData5[11238];
@(posedge clk);
#1;data_in = testData5[11239];
@(posedge clk);
#1;data_in = testData5[11240];
@(posedge clk);
#1;data_in = testData5[11241];
@(posedge clk);
#1;data_in = testData5[11242];
@(posedge clk);
#1;data_in = testData5[11243];
@(posedge clk);
#1;data_in = testData5[11244];
@(posedge clk);
#1;data_in = testData5[11245];
@(posedge clk);
#1;data_in = testData5[11246];
@(posedge clk);
#1;data_in = testData5[11247];
@(posedge clk);
#1;data_in = testData5[11248];
@(posedge clk);
#1;data_in = testData5[11249];
@(posedge clk);
#1;data_in = testData5[11250];
@(posedge clk);
#1;data_in = testData5[11251];
@(posedge clk);
#1;data_in = testData5[11252];
@(posedge clk);
#1;data_in = testData5[11253];
@(posedge clk);
#1;data_in = testData5[11254];
@(posedge clk);
#1;data_in = testData5[11255];
@(posedge clk);
#1;data_in = testData5[11256];
@(posedge clk);
#1;data_in = testData5[11257];
@(posedge clk);
#1;data_in = testData5[11258];
@(posedge clk);
#1;data_in = testData5[11259];
@(posedge clk);
#1;data_in = testData5[11260];
@(posedge clk);
#1;data_in = testData5[11261];
@(posedge clk);
#1;data_in = testData5[11262];
@(posedge clk);
#1;data_in = testData5[11263];
@(posedge clk);
#1;data_in = testData5[11264];
@(posedge clk);
#1;data_in = testData5[11265];
@(posedge clk);
#1;data_in = testData5[11266];
@(posedge clk);
#1;data_in = testData5[11267];
@(posedge clk);
#1;data_in = testData5[11268];
@(posedge clk);
#1;data_in = testData5[11269];
@(posedge clk);
#1;data_in = testData5[11270];
@(posedge clk);
#1;data_in = testData5[11271];
@(posedge clk);
#1;data_in = testData5[11272];
@(posedge clk);
#1;data_in = testData5[11273];
@(posedge clk);
#1;data_in = testData5[11274];
@(posedge clk);
#1;data_in = testData5[11275];
@(posedge clk);
#1;data_in = testData5[11276];
@(posedge clk);
#1;data_in = testData5[11277];
@(posedge clk);
#1;data_in = testData5[11278];
@(posedge clk);
#1;data_in = testData5[11279];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[11280]; 
@(posedge clk);
#1;data_in = testData5[11281];
@(posedge clk);
#1;data_in = testData5[11282];
@(posedge clk);
#1;data_in = testData5[11283];
@(posedge clk);
#1;data_in = testData5[11284];
@(posedge clk);
#1;data_in = testData5[11285];
@(posedge clk);
#1;data_in = testData5[11286];
@(posedge clk);
#1;data_in = testData5[11287];
@(posedge clk);
#1;data_in = testData5[11288];
@(posedge clk);
#1;data_in = testData5[11289];
@(posedge clk);
#1;data_in = testData5[11290];
@(posedge clk);
#1;data_in = testData5[11291];
@(posedge clk);
#1;data_in = testData5[11292];
@(posedge clk);
#1;data_in = testData5[11293];
@(posedge clk);
#1;data_in = testData5[11294];
@(posedge clk);
#1;data_in = testData5[11295];
@(posedge clk);
#1;data_in = testData5[11296];
@(posedge clk);
#1;data_in = testData5[11297];
@(posedge clk);
#1;data_in = testData5[11298];
@(posedge clk);
#1;data_in = testData5[11299];
@(posedge clk);
#1;data_in = testData5[11300];
@(posedge clk);
#1;data_in = testData5[11301];
@(posedge clk);
#1;data_in = testData5[11302];
@(posedge clk);
#1;data_in = testData5[11303];
@(posedge clk);
#1;data_in = testData5[11304];
@(posedge clk);
#1;data_in = testData5[11305];
@(posedge clk);
#1;data_in = testData5[11306];
@(posedge clk);
#1;data_in = testData5[11307];
@(posedge clk);
#1;data_in = testData5[11308];
@(posedge clk);
#1;data_in = testData5[11309];
@(posedge clk);
#1;data_in = testData5[11310];
@(posedge clk);
#1;data_in = testData5[11311];
@(posedge clk);
#1;data_in = testData5[11312];
@(posedge clk);
#1;data_in = testData5[11313];
@(posedge clk);
#1;data_in = testData5[11314];
@(posedge clk);
#1;data_in = testData5[11315];
@(posedge clk);
#1;data_in = testData5[11316];
@(posedge clk);
#1;data_in = testData5[11317];
@(posedge clk);
#1;data_in = testData5[11318];
@(posedge clk);
#1;data_in = testData5[11319];
@(posedge clk);
#1;data_in = testData5[11320];
@(posedge clk);
#1;data_in = testData5[11321];
@(posedge clk);
#1;data_in = testData5[11322];
@(posedge clk);
#1;data_in = testData5[11323];
@(posedge clk);
#1;data_in = testData5[11324];
@(posedge clk);
#1;data_in = testData5[11325];
@(posedge clk);
#1;data_in = testData5[11326];
@(posedge clk);
#1;data_in = testData5[11327];
@(posedge clk);
#1;data_in = testData5[11328];
@(posedge clk);
#1;data_in = testData5[11329];
@(posedge clk);
#1;data_in = testData5[11330];
@(posedge clk);
#1;data_in = testData5[11331];
@(posedge clk);
#1;data_in = testData5[11332];
@(posedge clk);
#1;data_in = testData5[11333];
@(posedge clk);
#1;data_in = testData5[11334];
@(posedge clk);
#1;data_in = testData5[11335];
@(posedge clk);
#1;data_in = testData5[11336];
@(posedge clk);
#1;data_in = testData5[11337];
@(posedge clk);
#1;data_in = testData5[11338];
@(posedge clk);
#1;data_in = testData5[11339];
@(posedge clk);
#1;data_in = testData5[11340];
@(posedge clk);
#1;data_in = testData5[11341];
@(posedge clk);
#1;data_in = testData5[11342];
@(posedge clk);
#1;data_in = testData5[11343];
@(posedge clk);
#1;data_in = testData5[11344];
@(posedge clk);
#1;data_in = testData5[11345];
@(posedge clk);
#1;data_in = testData5[11346];
@(posedge clk);
#1;data_in = testData5[11347];
@(posedge clk);
#1;data_in = testData5[11348];
@(posedge clk);
#1;data_in = testData5[11349];
@(posedge clk);
#1;data_in = testData5[11350];
@(posedge clk);
#1;data_in = testData5[11351];
@(posedge clk);
#1;data_in = testData5[11352];
@(posedge clk);
#1;data_in = testData5[11353];
@(posedge clk);
#1;data_in = testData5[11354];
@(posedge clk);
#1;data_in = testData5[11355];
@(posedge clk);
#1;data_in = testData5[11356];
@(posedge clk);
#1;data_in = testData5[11357];
@(posedge clk);
#1;data_in = testData5[11358];
@(posedge clk);
#1;data_in = testData5[11359];
@(posedge clk);
#1;data_in = testData5[11360];
@(posedge clk);
#1;data_in = testData5[11361];
@(posedge clk);
#1;data_in = testData5[11362];
@(posedge clk);
#1;data_in = testData5[11363];
@(posedge clk);
#1;data_in = testData5[11364];
@(posedge clk);
#1;data_in = testData5[11365];
@(posedge clk);
#1;data_in = testData5[11366];
@(posedge clk);
#1;data_in = testData5[11367];
@(posedge clk);
#1;data_in = testData5[11368];
@(posedge clk);
#1;data_in = testData5[11369];
@(posedge clk);
#1;data_in = testData5[11370];
@(posedge clk);
#1;data_in = testData5[11371];
@(posedge clk);
#1;data_in = testData5[11372];
@(posedge clk);
#1;data_in = testData5[11373];
@(posedge clk);
#1;data_in = testData5[11374];
@(posedge clk);
#1;data_in = testData5[11375];
@(posedge clk);
#1;data_in = testData5[11376];
@(posedge clk);
#1;data_in = testData5[11377];
@(posedge clk);
#1;data_in = testData5[11378];
@(posedge clk);
#1;data_in = testData5[11379];
@(posedge clk);
#1;data_in = testData5[11380];
@(posedge clk);
#1;data_in = testData5[11381];
@(posedge clk);
#1;data_in = testData5[11382];
@(posedge clk);
#1;data_in = testData5[11383];
@(posedge clk);
#1;data_in = testData5[11384];
@(posedge clk);
#1;data_in = testData5[11385];
@(posedge clk);
#1;data_in = testData5[11386];
@(posedge clk);
#1;data_in = testData5[11387];
@(posedge clk);
#1;data_in = testData5[11388];
@(posedge clk);
#1;data_in = testData5[11389];
@(posedge clk);
#1;data_in = testData5[11390];
@(posedge clk);
#1;data_in = testData5[11391];
@(posedge clk);
#1;data_in = testData5[11392];
@(posedge clk);
#1;data_in = testData5[11393];
@(posedge clk);
#1;data_in = testData5[11394];
@(posedge clk);
#1;data_in = testData5[11395];
@(posedge clk);
#1;data_in = testData5[11396];
@(posedge clk);
#1;data_in = testData5[11397];
@(posedge clk);
#1;data_in = testData5[11398];
@(posedge clk);
#1;data_in = testData5[11399];
@(posedge clk);
#1;data_in = testData5[11400];
@(posedge clk);
#1;data_in = testData5[11401];
@(posedge clk);
#1;data_in = testData5[11402];
@(posedge clk);
#1;data_in = testData5[11403];
@(posedge clk);
#1;data_in = testData5[11404];
@(posedge clk);
#1;data_in = testData5[11405];
@(posedge clk);
#1;data_in = testData5[11406];
@(posedge clk);
#1;data_in = testData5[11407];
@(posedge clk);
#1;data_in = testData5[11408];
@(posedge clk);
#1;data_in = testData5[11409];
@(posedge clk);
#1;data_in = testData5[11410];
@(posedge clk);
#1;data_in = testData5[11411];
@(posedge clk);
#1;data_in = testData5[11412];
@(posedge clk);
#1;data_in = testData5[11413];
@(posedge clk);
#1;data_in = testData5[11414];
@(posedge clk);
#1;data_in = testData5[11415];
@(posedge clk);
#1;data_in = testData5[11416];
@(posedge clk);
#1;data_in = testData5[11417];
@(posedge clk);
#1;data_in = testData5[11418];
@(posedge clk);
#1;data_in = testData5[11419];
@(posedge clk);
#1;data_in = testData5[11420];
@(posedge clk);
#1;data_in = testData5[11421];
@(posedge clk);
#1;data_in = testData5[11422];
@(posedge clk);
#1;data_in = testData5[11423];
@(posedge clk);
#1;data_in = testData5[11424];
@(posedge clk);
#1;data_in = testData5[11425];
@(posedge clk);
#1;data_in = testData5[11426];
@(posedge clk);
#1;data_in = testData5[11427];
@(posedge clk);
#1;data_in = testData5[11428];
@(posedge clk);
#1;data_in = testData5[11429];
@(posedge clk);
#1;data_in = testData5[11430];
@(posedge clk);
#1;data_in = testData5[11431];
@(posedge clk);
#1;data_in = testData5[11432];
@(posedge clk);
#1;data_in = testData5[11433];
@(posedge clk);
#1;data_in = testData5[11434];
@(posedge clk);
#1;data_in = testData5[11435];
@(posedge clk);
#1;data_in = testData5[11436];
@(posedge clk);
#1;data_in = testData5[11437];
@(posedge clk);
#1;data_in = testData5[11438];
@(posedge clk);
#1;data_in = testData5[11439];
@(posedge clk);
#1;data_in = testData5[11440];
@(posedge clk);
#1;data_in = testData5[11441];
@(posedge clk);
#1;data_in = testData5[11442];
@(posedge clk);
#1;data_in = testData5[11443];
@(posedge clk);
#1;data_in = testData5[11444];
@(posedge clk);
#1;data_in = testData5[11445];
@(posedge clk);
#1;data_in = testData5[11446];
@(posedge clk);
#1;data_in = testData5[11447];
@(posedge clk);
#1;data_in = testData5[11448];
@(posedge clk);
#1;data_in = testData5[11449];
@(posedge clk);
#1;data_in = testData5[11450];
@(posedge clk);
#1;data_in = testData5[11451];
@(posedge clk);
#1;data_in = testData5[11452];
@(posedge clk);
#1;data_in = testData5[11453];
@(posedge clk);
#1;data_in = testData5[11454];
@(posedge clk);
#1;data_in = testData5[11455];
@(posedge clk);
#1;data_in = testData5[11456];
@(posedge clk);
#1;data_in = testData5[11457];
@(posedge clk);
#1;data_in = testData5[11458];
@(posedge clk);
#1;data_in = testData5[11459];
@(posedge clk);
#1;data_in = testData5[11460];
@(posedge clk);
#1;data_in = testData5[11461];
@(posedge clk);
#1;data_in = testData5[11462];
@(posedge clk);
#1;data_in = testData5[11463];
@(posedge clk);
#1;data_in = testData5[11464];
@(posedge clk);
#1;data_in = testData5[11465];
@(posedge clk);
#1;data_in = testData5[11466];
@(posedge clk);
#1;data_in = testData5[11467];
@(posedge clk);
#1;data_in = testData5[11468];
@(posedge clk);
#1;data_in = testData5[11469];
@(posedge clk);
#1;data_in = testData5[11470];
@(posedge clk);
#1;data_in = testData5[11471];
@(posedge clk);
#1;data_in = testData5[11472];
@(posedge clk);
#1;data_in = testData5[11473];
@(posedge clk);
#1;data_in = testData5[11474];
@(posedge clk);
#1;data_in = testData5[11475];
@(posedge clk);
#1;data_in = testData5[11476];
@(posedge clk);
#1;data_in = testData5[11477];
@(posedge clk);
#1;data_in = testData5[11478];
@(posedge clk);
#1;data_in = testData5[11479];
@(posedge clk);
#1;data_in = testData5[11480];
@(posedge clk);
#1;data_in = testData5[11481];
@(posedge clk);
#1;data_in = testData5[11482];
@(posedge clk);
#1;data_in = testData5[11483];
@(posedge clk);
#1;data_in = testData5[11484];
@(posedge clk);
#1;data_in = testData5[11485];
@(posedge clk);
#1;data_in = testData5[11486];
@(posedge clk);
#1;data_in = testData5[11487];
@(posedge clk);
#1;data_in = testData5[11488];
@(posedge clk);
#1;data_in = testData5[11489];
@(posedge clk);
#1;data_in = testData5[11490];
@(posedge clk);
#1;data_in = testData5[11491];
@(posedge clk);
#1;data_in = testData5[11492];
@(posedge clk);
#1;data_in = testData5[11493];
@(posedge clk);
#1;data_in = testData5[11494];
@(posedge clk);
#1;data_in = testData5[11495];
@(posedge clk);
#1;data_in = testData5[11496];
@(posedge clk);
#1;data_in = testData5[11497];
@(posedge clk);
#1;data_in = testData5[11498];
@(posedge clk);
#1;data_in = testData5[11499];
@(posedge clk);
#1;data_in = testData5[11500];
@(posedge clk);
#1;data_in = testData5[11501];
@(posedge clk);
#1;data_in = testData5[11502];
@(posedge clk);
#1;data_in = testData5[11503];
@(posedge clk);
#1;data_in = testData5[11504];
@(posedge clk);
#1;data_in = testData5[11505];
@(posedge clk);
#1;data_in = testData5[11506];
@(posedge clk);
#1;data_in = testData5[11507];
@(posedge clk);
#1;data_in = testData5[11508];
@(posedge clk);
#1;data_in = testData5[11509];
@(posedge clk);
#1;data_in = testData5[11510];
@(posedge clk);
#1;data_in = testData5[11511];
@(posedge clk);
#1;data_in = testData5[11512];
@(posedge clk);
#1;data_in = testData5[11513];
@(posedge clk);
#1;data_in = testData5[11514];
@(posedge clk);
#1;data_in = testData5[11515];
@(posedge clk);
#1;data_in = testData5[11516];
@(posedge clk);
#1;data_in = testData5[11517];
@(posedge clk);
#1;data_in = testData5[11518];
@(posedge clk);
#1;data_in = testData5[11519];
@(posedge clk);
#1;data_in = testData5[11520];
@(posedge clk);
#1;data_in = testData5[11521];
@(posedge clk);
#1;data_in = testData5[11522];
@(posedge clk);
#1;data_in = testData5[11523];
@(posedge clk);
#1;data_in = testData5[11524];
@(posedge clk);
#1;data_in = testData5[11525];
@(posedge clk);
#1;data_in = testData5[11526];
@(posedge clk);
#1;data_in = testData5[11527];
@(posedge clk);
#1;data_in = testData5[11528];
@(posedge clk);
#1;data_in = testData5[11529];
@(posedge clk);
#1;data_in = testData5[11530];
@(posedge clk);
#1;data_in = testData5[11531];
@(posedge clk);
#1;data_in = testData5[11532];
@(posedge clk);
#1;data_in = testData5[11533];
@(posedge clk);
#1;data_in = testData5[11534];
@(posedge clk);
#1;data_in = testData5[11535];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[11536]; 
@(posedge clk);
#1;data_in = testData5[11537];
@(posedge clk);
#1;data_in = testData5[11538];
@(posedge clk);
#1;data_in = testData5[11539];
@(posedge clk);
#1;data_in = testData5[11540];
@(posedge clk);
#1;data_in = testData5[11541];
@(posedge clk);
#1;data_in = testData5[11542];
@(posedge clk);
#1;data_in = testData5[11543];
@(posedge clk);
#1;data_in = testData5[11544];
@(posedge clk);
#1;data_in = testData5[11545];
@(posedge clk);
#1;data_in = testData5[11546];
@(posedge clk);
#1;data_in = testData5[11547];
@(posedge clk);
#1;data_in = testData5[11548];
@(posedge clk);
#1;data_in = testData5[11549];
@(posedge clk);
#1;data_in = testData5[11550];
@(posedge clk);
#1;data_in = testData5[11551];
@(posedge clk);
#1;data_in = testData5[11552];
@(posedge clk);
#1;data_in = testData5[11553];
@(posedge clk);
#1;data_in = testData5[11554];
@(posedge clk);
#1;data_in = testData5[11555];
@(posedge clk);
#1;data_in = testData5[11556];
@(posedge clk);
#1;data_in = testData5[11557];
@(posedge clk);
#1;data_in = testData5[11558];
@(posedge clk);
#1;data_in = testData5[11559];
@(posedge clk);
#1;data_in = testData5[11560];
@(posedge clk);
#1;data_in = testData5[11561];
@(posedge clk);
#1;data_in = testData5[11562];
@(posedge clk);
#1;data_in = testData5[11563];
@(posedge clk);
#1;data_in = testData5[11564];
@(posedge clk);
#1;data_in = testData5[11565];
@(posedge clk);
#1;data_in = testData5[11566];
@(posedge clk);
#1;data_in = testData5[11567];
@(posedge clk);
#1;data_in = testData5[11568];
@(posedge clk);
#1;data_in = testData5[11569];
@(posedge clk);
#1;data_in = testData5[11570];
@(posedge clk);
#1;data_in = testData5[11571];
@(posedge clk);
#1;data_in = testData5[11572];
@(posedge clk);
#1;data_in = testData5[11573];
@(posedge clk);
#1;data_in = testData5[11574];
@(posedge clk);
#1;data_in = testData5[11575];
@(posedge clk);
#1;data_in = testData5[11576];
@(posedge clk);
#1;data_in = testData5[11577];
@(posedge clk);
#1;data_in = testData5[11578];
@(posedge clk);
#1;data_in = testData5[11579];
@(posedge clk);
#1;data_in = testData5[11580];
@(posedge clk);
#1;data_in = testData5[11581];
@(posedge clk);
#1;data_in = testData5[11582];
@(posedge clk);
#1;data_in = testData5[11583];
@(posedge clk);
#1;data_in = testData5[11584];
@(posedge clk);
#1;data_in = testData5[11585];
@(posedge clk);
#1;data_in = testData5[11586];
@(posedge clk);
#1;data_in = testData5[11587];
@(posedge clk);
#1;data_in = testData5[11588];
@(posedge clk);
#1;data_in = testData5[11589];
@(posedge clk);
#1;data_in = testData5[11590];
@(posedge clk);
#1;data_in = testData5[11591];
@(posedge clk);
#1;data_in = testData5[11592];
@(posedge clk);
#1;data_in = testData5[11593];
@(posedge clk);
#1;data_in = testData5[11594];
@(posedge clk);
#1;data_in = testData5[11595];
@(posedge clk);
#1;data_in = testData5[11596];
@(posedge clk);
#1;data_in = testData5[11597];
@(posedge clk);
#1;data_in = testData5[11598];
@(posedge clk);
#1;data_in = testData5[11599];
@(posedge clk);
#1;data_in = testData5[11600];
@(posedge clk);
#1;data_in = testData5[11601];
@(posedge clk);
#1;data_in = testData5[11602];
@(posedge clk);
#1;data_in = testData5[11603];
@(posedge clk);
#1;data_in = testData5[11604];
@(posedge clk);
#1;data_in = testData5[11605];
@(posedge clk);
#1;data_in = testData5[11606];
@(posedge clk);
#1;data_in = testData5[11607];
@(posedge clk);
#1;data_in = testData5[11608];
@(posedge clk);
#1;data_in = testData5[11609];
@(posedge clk);
#1;data_in = testData5[11610];
@(posedge clk);
#1;data_in = testData5[11611];
@(posedge clk);
#1;data_in = testData5[11612];
@(posedge clk);
#1;data_in = testData5[11613];
@(posedge clk);
#1;data_in = testData5[11614];
@(posedge clk);
#1;data_in = testData5[11615];
@(posedge clk);
#1;data_in = testData5[11616];
@(posedge clk);
#1;data_in = testData5[11617];
@(posedge clk);
#1;data_in = testData5[11618];
@(posedge clk);
#1;data_in = testData5[11619];
@(posedge clk);
#1;data_in = testData5[11620];
@(posedge clk);
#1;data_in = testData5[11621];
@(posedge clk);
#1;data_in = testData5[11622];
@(posedge clk);
#1;data_in = testData5[11623];
@(posedge clk);
#1;data_in = testData5[11624];
@(posedge clk);
#1;data_in = testData5[11625];
@(posedge clk);
#1;data_in = testData5[11626];
@(posedge clk);
#1;data_in = testData5[11627];
@(posedge clk);
#1;data_in = testData5[11628];
@(posedge clk);
#1;data_in = testData5[11629];
@(posedge clk);
#1;data_in = testData5[11630];
@(posedge clk);
#1;data_in = testData5[11631];
@(posedge clk);
#1;data_in = testData5[11632];
@(posedge clk);
#1;data_in = testData5[11633];
@(posedge clk);
#1;data_in = testData5[11634];
@(posedge clk);
#1;data_in = testData5[11635];
@(posedge clk);
#1;data_in = testData5[11636];
@(posedge clk);
#1;data_in = testData5[11637];
@(posedge clk);
#1;data_in = testData5[11638];
@(posedge clk);
#1;data_in = testData5[11639];
@(posedge clk);
#1;data_in = testData5[11640];
@(posedge clk);
#1;data_in = testData5[11641];
@(posedge clk);
#1;data_in = testData5[11642];
@(posedge clk);
#1;data_in = testData5[11643];
@(posedge clk);
#1;data_in = testData5[11644];
@(posedge clk);
#1;data_in = testData5[11645];
@(posedge clk);
#1;data_in = testData5[11646];
@(posedge clk);
#1;data_in = testData5[11647];
@(posedge clk);
#1;data_in = testData5[11648];
@(posedge clk);
#1;data_in = testData5[11649];
@(posedge clk);
#1;data_in = testData5[11650];
@(posedge clk);
#1;data_in = testData5[11651];
@(posedge clk);
#1;data_in = testData5[11652];
@(posedge clk);
#1;data_in = testData5[11653];
@(posedge clk);
#1;data_in = testData5[11654];
@(posedge clk);
#1;data_in = testData5[11655];
@(posedge clk);
#1;data_in = testData5[11656];
@(posedge clk);
#1;data_in = testData5[11657];
@(posedge clk);
#1;data_in = testData5[11658];
@(posedge clk);
#1;data_in = testData5[11659];
@(posedge clk);
#1;data_in = testData5[11660];
@(posedge clk);
#1;data_in = testData5[11661];
@(posedge clk);
#1;data_in = testData5[11662];
@(posedge clk);
#1;data_in = testData5[11663];
@(posedge clk);
#1;data_in = testData5[11664];
@(posedge clk);
#1;data_in = testData5[11665];
@(posedge clk);
#1;data_in = testData5[11666];
@(posedge clk);
#1;data_in = testData5[11667];
@(posedge clk);
#1;data_in = testData5[11668];
@(posedge clk);
#1;data_in = testData5[11669];
@(posedge clk);
#1;data_in = testData5[11670];
@(posedge clk);
#1;data_in = testData5[11671];
@(posedge clk);
#1;data_in = testData5[11672];
@(posedge clk);
#1;data_in = testData5[11673];
@(posedge clk);
#1;data_in = testData5[11674];
@(posedge clk);
#1;data_in = testData5[11675];
@(posedge clk);
#1;data_in = testData5[11676];
@(posedge clk);
#1;data_in = testData5[11677];
@(posedge clk);
#1;data_in = testData5[11678];
@(posedge clk);
#1;data_in = testData5[11679];
@(posedge clk);
#1;data_in = testData5[11680];
@(posedge clk);
#1;data_in = testData5[11681];
@(posedge clk);
#1;data_in = testData5[11682];
@(posedge clk);
#1;data_in = testData5[11683];
@(posedge clk);
#1;data_in = testData5[11684];
@(posedge clk);
#1;data_in = testData5[11685];
@(posedge clk);
#1;data_in = testData5[11686];
@(posedge clk);
#1;data_in = testData5[11687];
@(posedge clk);
#1;data_in = testData5[11688];
@(posedge clk);
#1;data_in = testData5[11689];
@(posedge clk);
#1;data_in = testData5[11690];
@(posedge clk);
#1;data_in = testData5[11691];
@(posedge clk);
#1;data_in = testData5[11692];
@(posedge clk);
#1;data_in = testData5[11693];
@(posedge clk);
#1;data_in = testData5[11694];
@(posedge clk);
#1;data_in = testData5[11695];
@(posedge clk);
#1;data_in = testData5[11696];
@(posedge clk);
#1;data_in = testData5[11697];
@(posedge clk);
#1;data_in = testData5[11698];
@(posedge clk);
#1;data_in = testData5[11699];
@(posedge clk);
#1;data_in = testData5[11700];
@(posedge clk);
#1;data_in = testData5[11701];
@(posedge clk);
#1;data_in = testData5[11702];
@(posedge clk);
#1;data_in = testData5[11703];
@(posedge clk);
#1;data_in = testData5[11704];
@(posedge clk);
#1;data_in = testData5[11705];
@(posedge clk);
#1;data_in = testData5[11706];
@(posedge clk);
#1;data_in = testData5[11707];
@(posedge clk);
#1;data_in = testData5[11708];
@(posedge clk);
#1;data_in = testData5[11709];
@(posedge clk);
#1;data_in = testData5[11710];
@(posedge clk);
#1;data_in = testData5[11711];
@(posedge clk);
#1;data_in = testData5[11712];
@(posedge clk);
#1;data_in = testData5[11713];
@(posedge clk);
#1;data_in = testData5[11714];
@(posedge clk);
#1;data_in = testData5[11715];
@(posedge clk);
#1;data_in = testData5[11716];
@(posedge clk);
#1;data_in = testData5[11717];
@(posedge clk);
#1;data_in = testData5[11718];
@(posedge clk);
#1;data_in = testData5[11719];
@(posedge clk);
#1;data_in = testData5[11720];
@(posedge clk);
#1;data_in = testData5[11721];
@(posedge clk);
#1;data_in = testData5[11722];
@(posedge clk);
#1;data_in = testData5[11723];
@(posedge clk);
#1;data_in = testData5[11724];
@(posedge clk);
#1;data_in = testData5[11725];
@(posedge clk);
#1;data_in = testData5[11726];
@(posedge clk);
#1;data_in = testData5[11727];
@(posedge clk);
#1;data_in = testData5[11728];
@(posedge clk);
#1;data_in = testData5[11729];
@(posedge clk);
#1;data_in = testData5[11730];
@(posedge clk);
#1;data_in = testData5[11731];
@(posedge clk);
#1;data_in = testData5[11732];
@(posedge clk);
#1;data_in = testData5[11733];
@(posedge clk);
#1;data_in = testData5[11734];
@(posedge clk);
#1;data_in = testData5[11735];
@(posedge clk);
#1;data_in = testData5[11736];
@(posedge clk);
#1;data_in = testData5[11737];
@(posedge clk);
#1;data_in = testData5[11738];
@(posedge clk);
#1;data_in = testData5[11739];
@(posedge clk);
#1;data_in = testData5[11740];
@(posedge clk);
#1;data_in = testData5[11741];
@(posedge clk);
#1;data_in = testData5[11742];
@(posedge clk);
#1;data_in = testData5[11743];
@(posedge clk);
#1;data_in = testData5[11744];
@(posedge clk);
#1;data_in = testData5[11745];
@(posedge clk);
#1;data_in = testData5[11746];
@(posedge clk);
#1;data_in = testData5[11747];
@(posedge clk);
#1;data_in = testData5[11748];
@(posedge clk);
#1;data_in = testData5[11749];
@(posedge clk);
#1;data_in = testData5[11750];
@(posedge clk);
#1;data_in = testData5[11751];
@(posedge clk);
#1;data_in = testData5[11752];
@(posedge clk);
#1;data_in = testData5[11753];
@(posedge clk);
#1;data_in = testData5[11754];
@(posedge clk);
#1;data_in = testData5[11755];
@(posedge clk);
#1;data_in = testData5[11756];
@(posedge clk);
#1;data_in = testData5[11757];
@(posedge clk);
#1;data_in = testData5[11758];
@(posedge clk);
#1;data_in = testData5[11759];
@(posedge clk);
#1;data_in = testData5[11760];
@(posedge clk);
#1;data_in = testData5[11761];
@(posedge clk);
#1;data_in = testData5[11762];
@(posedge clk);
#1;data_in = testData5[11763];
@(posedge clk);
#1;data_in = testData5[11764];
@(posedge clk);
#1;data_in = testData5[11765];
@(posedge clk);
#1;data_in = testData5[11766];
@(posedge clk);
#1;data_in = testData5[11767];
@(posedge clk);
#1;data_in = testData5[11768];
@(posedge clk);
#1;data_in = testData5[11769];
@(posedge clk);
#1;data_in = testData5[11770];
@(posedge clk);
#1;data_in = testData5[11771];
@(posedge clk);
#1;data_in = testData5[11772];
@(posedge clk);
#1;data_in = testData5[11773];
@(posedge clk);
#1;data_in = testData5[11774];
@(posedge clk);
#1;data_in = testData5[11775];
@(posedge clk);
#1;data_in = testData5[11776];
@(posedge clk);
#1;data_in = testData5[11777];
@(posedge clk);
#1;data_in = testData5[11778];
@(posedge clk);
#1;data_in = testData5[11779];
@(posedge clk);
#1;data_in = testData5[11780];
@(posedge clk);
#1;data_in = testData5[11781];
@(posedge clk);
#1;data_in = testData5[11782];
@(posedge clk);
#1;data_in = testData5[11783];
@(posedge clk);
#1;data_in = testData5[11784];
@(posedge clk);
#1;data_in = testData5[11785];
@(posedge clk);
#1;data_in = testData5[11786];
@(posedge clk);
#1;data_in = testData5[11787];
@(posedge clk);
#1;data_in = testData5[11788];
@(posedge clk);
#1;data_in = testData5[11789];
@(posedge clk);
#1;data_in = testData5[11790];
@(posedge clk);
#1;data_in = testData5[11791];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[11792]; 
@(posedge clk);
#1;data_in = testData5[11793];
@(posedge clk);
#1;data_in = testData5[11794];
@(posedge clk);
#1;data_in = testData5[11795];
@(posedge clk);
#1;data_in = testData5[11796];
@(posedge clk);
#1;data_in = testData5[11797];
@(posedge clk);
#1;data_in = testData5[11798];
@(posedge clk);
#1;data_in = testData5[11799];
@(posedge clk);
#1;data_in = testData5[11800];
@(posedge clk);
#1;data_in = testData5[11801];
@(posedge clk);
#1;data_in = testData5[11802];
@(posedge clk);
#1;data_in = testData5[11803];
@(posedge clk);
#1;data_in = testData5[11804];
@(posedge clk);
#1;data_in = testData5[11805];
@(posedge clk);
#1;data_in = testData5[11806];
@(posedge clk);
#1;data_in = testData5[11807];
@(posedge clk);
#1;data_in = testData5[11808];
@(posedge clk);
#1;data_in = testData5[11809];
@(posedge clk);
#1;data_in = testData5[11810];
@(posedge clk);
#1;data_in = testData5[11811];
@(posedge clk);
#1;data_in = testData5[11812];
@(posedge clk);
#1;data_in = testData5[11813];
@(posedge clk);
#1;data_in = testData5[11814];
@(posedge clk);
#1;data_in = testData5[11815];
@(posedge clk);
#1;data_in = testData5[11816];
@(posedge clk);
#1;data_in = testData5[11817];
@(posedge clk);
#1;data_in = testData5[11818];
@(posedge clk);
#1;data_in = testData5[11819];
@(posedge clk);
#1;data_in = testData5[11820];
@(posedge clk);
#1;data_in = testData5[11821];
@(posedge clk);
#1;data_in = testData5[11822];
@(posedge clk);
#1;data_in = testData5[11823];
@(posedge clk);
#1;data_in = testData5[11824];
@(posedge clk);
#1;data_in = testData5[11825];
@(posedge clk);
#1;data_in = testData5[11826];
@(posedge clk);
#1;data_in = testData5[11827];
@(posedge clk);
#1;data_in = testData5[11828];
@(posedge clk);
#1;data_in = testData5[11829];
@(posedge clk);
#1;data_in = testData5[11830];
@(posedge clk);
#1;data_in = testData5[11831];
@(posedge clk);
#1;data_in = testData5[11832];
@(posedge clk);
#1;data_in = testData5[11833];
@(posedge clk);
#1;data_in = testData5[11834];
@(posedge clk);
#1;data_in = testData5[11835];
@(posedge clk);
#1;data_in = testData5[11836];
@(posedge clk);
#1;data_in = testData5[11837];
@(posedge clk);
#1;data_in = testData5[11838];
@(posedge clk);
#1;data_in = testData5[11839];
@(posedge clk);
#1;data_in = testData5[11840];
@(posedge clk);
#1;data_in = testData5[11841];
@(posedge clk);
#1;data_in = testData5[11842];
@(posedge clk);
#1;data_in = testData5[11843];
@(posedge clk);
#1;data_in = testData5[11844];
@(posedge clk);
#1;data_in = testData5[11845];
@(posedge clk);
#1;data_in = testData5[11846];
@(posedge clk);
#1;data_in = testData5[11847];
@(posedge clk);
#1;data_in = testData5[11848];
@(posedge clk);
#1;data_in = testData5[11849];
@(posedge clk);
#1;data_in = testData5[11850];
@(posedge clk);
#1;data_in = testData5[11851];
@(posedge clk);
#1;data_in = testData5[11852];
@(posedge clk);
#1;data_in = testData5[11853];
@(posedge clk);
#1;data_in = testData5[11854];
@(posedge clk);
#1;data_in = testData5[11855];
@(posedge clk);
#1;data_in = testData5[11856];
@(posedge clk);
#1;data_in = testData5[11857];
@(posedge clk);
#1;data_in = testData5[11858];
@(posedge clk);
#1;data_in = testData5[11859];
@(posedge clk);
#1;data_in = testData5[11860];
@(posedge clk);
#1;data_in = testData5[11861];
@(posedge clk);
#1;data_in = testData5[11862];
@(posedge clk);
#1;data_in = testData5[11863];
@(posedge clk);
#1;data_in = testData5[11864];
@(posedge clk);
#1;data_in = testData5[11865];
@(posedge clk);
#1;data_in = testData5[11866];
@(posedge clk);
#1;data_in = testData5[11867];
@(posedge clk);
#1;data_in = testData5[11868];
@(posedge clk);
#1;data_in = testData5[11869];
@(posedge clk);
#1;data_in = testData5[11870];
@(posedge clk);
#1;data_in = testData5[11871];
@(posedge clk);
#1;data_in = testData5[11872];
@(posedge clk);
#1;data_in = testData5[11873];
@(posedge clk);
#1;data_in = testData5[11874];
@(posedge clk);
#1;data_in = testData5[11875];
@(posedge clk);
#1;data_in = testData5[11876];
@(posedge clk);
#1;data_in = testData5[11877];
@(posedge clk);
#1;data_in = testData5[11878];
@(posedge clk);
#1;data_in = testData5[11879];
@(posedge clk);
#1;data_in = testData5[11880];
@(posedge clk);
#1;data_in = testData5[11881];
@(posedge clk);
#1;data_in = testData5[11882];
@(posedge clk);
#1;data_in = testData5[11883];
@(posedge clk);
#1;data_in = testData5[11884];
@(posedge clk);
#1;data_in = testData5[11885];
@(posedge clk);
#1;data_in = testData5[11886];
@(posedge clk);
#1;data_in = testData5[11887];
@(posedge clk);
#1;data_in = testData5[11888];
@(posedge clk);
#1;data_in = testData5[11889];
@(posedge clk);
#1;data_in = testData5[11890];
@(posedge clk);
#1;data_in = testData5[11891];
@(posedge clk);
#1;data_in = testData5[11892];
@(posedge clk);
#1;data_in = testData5[11893];
@(posedge clk);
#1;data_in = testData5[11894];
@(posedge clk);
#1;data_in = testData5[11895];
@(posedge clk);
#1;data_in = testData5[11896];
@(posedge clk);
#1;data_in = testData5[11897];
@(posedge clk);
#1;data_in = testData5[11898];
@(posedge clk);
#1;data_in = testData5[11899];
@(posedge clk);
#1;data_in = testData5[11900];
@(posedge clk);
#1;data_in = testData5[11901];
@(posedge clk);
#1;data_in = testData5[11902];
@(posedge clk);
#1;data_in = testData5[11903];
@(posedge clk);
#1;data_in = testData5[11904];
@(posedge clk);
#1;data_in = testData5[11905];
@(posedge clk);
#1;data_in = testData5[11906];
@(posedge clk);
#1;data_in = testData5[11907];
@(posedge clk);
#1;data_in = testData5[11908];
@(posedge clk);
#1;data_in = testData5[11909];
@(posedge clk);
#1;data_in = testData5[11910];
@(posedge clk);
#1;data_in = testData5[11911];
@(posedge clk);
#1;data_in = testData5[11912];
@(posedge clk);
#1;data_in = testData5[11913];
@(posedge clk);
#1;data_in = testData5[11914];
@(posedge clk);
#1;data_in = testData5[11915];
@(posedge clk);
#1;data_in = testData5[11916];
@(posedge clk);
#1;data_in = testData5[11917];
@(posedge clk);
#1;data_in = testData5[11918];
@(posedge clk);
#1;data_in = testData5[11919];
@(posedge clk);
#1;data_in = testData5[11920];
@(posedge clk);
#1;data_in = testData5[11921];
@(posedge clk);
#1;data_in = testData5[11922];
@(posedge clk);
#1;data_in = testData5[11923];
@(posedge clk);
#1;data_in = testData5[11924];
@(posedge clk);
#1;data_in = testData5[11925];
@(posedge clk);
#1;data_in = testData5[11926];
@(posedge clk);
#1;data_in = testData5[11927];
@(posedge clk);
#1;data_in = testData5[11928];
@(posedge clk);
#1;data_in = testData5[11929];
@(posedge clk);
#1;data_in = testData5[11930];
@(posedge clk);
#1;data_in = testData5[11931];
@(posedge clk);
#1;data_in = testData5[11932];
@(posedge clk);
#1;data_in = testData5[11933];
@(posedge clk);
#1;data_in = testData5[11934];
@(posedge clk);
#1;data_in = testData5[11935];
@(posedge clk);
#1;data_in = testData5[11936];
@(posedge clk);
#1;data_in = testData5[11937];
@(posedge clk);
#1;data_in = testData5[11938];
@(posedge clk);
#1;data_in = testData5[11939];
@(posedge clk);
#1;data_in = testData5[11940];
@(posedge clk);
#1;data_in = testData5[11941];
@(posedge clk);
#1;data_in = testData5[11942];
@(posedge clk);
#1;data_in = testData5[11943];
@(posedge clk);
#1;data_in = testData5[11944];
@(posedge clk);
#1;data_in = testData5[11945];
@(posedge clk);
#1;data_in = testData5[11946];
@(posedge clk);
#1;data_in = testData5[11947];
@(posedge clk);
#1;data_in = testData5[11948];
@(posedge clk);
#1;data_in = testData5[11949];
@(posedge clk);
#1;data_in = testData5[11950];
@(posedge clk);
#1;data_in = testData5[11951];
@(posedge clk);
#1;data_in = testData5[11952];
@(posedge clk);
#1;data_in = testData5[11953];
@(posedge clk);
#1;data_in = testData5[11954];
@(posedge clk);
#1;data_in = testData5[11955];
@(posedge clk);
#1;data_in = testData5[11956];
@(posedge clk);
#1;data_in = testData5[11957];
@(posedge clk);
#1;data_in = testData5[11958];
@(posedge clk);
#1;data_in = testData5[11959];
@(posedge clk);
#1;data_in = testData5[11960];
@(posedge clk);
#1;data_in = testData5[11961];
@(posedge clk);
#1;data_in = testData5[11962];
@(posedge clk);
#1;data_in = testData5[11963];
@(posedge clk);
#1;data_in = testData5[11964];
@(posedge clk);
#1;data_in = testData5[11965];
@(posedge clk);
#1;data_in = testData5[11966];
@(posedge clk);
#1;data_in = testData5[11967];
@(posedge clk);
#1;data_in = testData5[11968];
@(posedge clk);
#1;data_in = testData5[11969];
@(posedge clk);
#1;data_in = testData5[11970];
@(posedge clk);
#1;data_in = testData5[11971];
@(posedge clk);
#1;data_in = testData5[11972];
@(posedge clk);
#1;data_in = testData5[11973];
@(posedge clk);
#1;data_in = testData5[11974];
@(posedge clk);
#1;data_in = testData5[11975];
@(posedge clk);
#1;data_in = testData5[11976];
@(posedge clk);
#1;data_in = testData5[11977];
@(posedge clk);
#1;data_in = testData5[11978];
@(posedge clk);
#1;data_in = testData5[11979];
@(posedge clk);
#1;data_in = testData5[11980];
@(posedge clk);
#1;data_in = testData5[11981];
@(posedge clk);
#1;data_in = testData5[11982];
@(posedge clk);
#1;data_in = testData5[11983];
@(posedge clk);
#1;data_in = testData5[11984];
@(posedge clk);
#1;data_in = testData5[11985];
@(posedge clk);
#1;data_in = testData5[11986];
@(posedge clk);
#1;data_in = testData5[11987];
@(posedge clk);
#1;data_in = testData5[11988];
@(posedge clk);
#1;data_in = testData5[11989];
@(posedge clk);
#1;data_in = testData5[11990];
@(posedge clk);
#1;data_in = testData5[11991];
@(posedge clk);
#1;data_in = testData5[11992];
@(posedge clk);
#1;data_in = testData5[11993];
@(posedge clk);
#1;data_in = testData5[11994];
@(posedge clk);
#1;data_in = testData5[11995];
@(posedge clk);
#1;data_in = testData5[11996];
@(posedge clk);
#1;data_in = testData5[11997];
@(posedge clk);
#1;data_in = testData5[11998];
@(posedge clk);
#1;data_in = testData5[11999];
@(posedge clk);
#1;data_in = testData5[12000];
@(posedge clk);
#1;data_in = testData5[12001];
@(posedge clk);
#1;data_in = testData5[12002];
@(posedge clk);
#1;data_in = testData5[12003];
@(posedge clk);
#1;data_in = testData5[12004];
@(posedge clk);
#1;data_in = testData5[12005];
@(posedge clk);
#1;data_in = testData5[12006];
@(posedge clk);
#1;data_in = testData5[12007];
@(posedge clk);
#1;data_in = testData5[12008];
@(posedge clk);
#1;data_in = testData5[12009];
@(posedge clk);
#1;data_in = testData5[12010];
@(posedge clk);
#1;data_in = testData5[12011];
@(posedge clk);
#1;data_in = testData5[12012];
@(posedge clk);
#1;data_in = testData5[12013];
@(posedge clk);
#1;data_in = testData5[12014];
@(posedge clk);
#1;data_in = testData5[12015];
@(posedge clk);
#1;data_in = testData5[12016];
@(posedge clk);
#1;data_in = testData5[12017];
@(posedge clk);
#1;data_in = testData5[12018];
@(posedge clk);
#1;data_in = testData5[12019];
@(posedge clk);
#1;data_in = testData5[12020];
@(posedge clk);
#1;data_in = testData5[12021];
@(posedge clk);
#1;data_in = testData5[12022];
@(posedge clk);
#1;data_in = testData5[12023];
@(posedge clk);
#1;data_in = testData5[12024];
@(posedge clk);
#1;data_in = testData5[12025];
@(posedge clk);
#1;data_in = testData5[12026];
@(posedge clk);
#1;data_in = testData5[12027];
@(posedge clk);
#1;data_in = testData5[12028];
@(posedge clk);
#1;data_in = testData5[12029];
@(posedge clk);
#1;data_in = testData5[12030];
@(posedge clk);
#1;data_in = testData5[12031];
@(posedge clk);
#1;data_in = testData5[12032];
@(posedge clk);
#1;data_in = testData5[12033];
@(posedge clk);
#1;data_in = testData5[12034];
@(posedge clk);
#1;data_in = testData5[12035];
@(posedge clk);
#1;data_in = testData5[12036];
@(posedge clk);
#1;data_in = testData5[12037];
@(posedge clk);
#1;data_in = testData5[12038];
@(posedge clk);
#1;data_in = testData5[12039];
@(posedge clk);
#1;data_in = testData5[12040];
@(posedge clk);
#1;data_in = testData5[12041];
@(posedge clk);
#1;data_in = testData5[12042];
@(posedge clk);
#1;data_in = testData5[12043];
@(posedge clk);
#1;data_in = testData5[12044];
@(posedge clk);
#1;data_in = testData5[12045];
@(posedge clk);
#1;data_in = testData5[12046];
@(posedge clk);
#1;data_in = testData5[12047];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[12048]; 
@(posedge clk);
#1;data_in = testData5[12049];
@(posedge clk);
#1;data_in = testData5[12050];
@(posedge clk);
#1;data_in = testData5[12051];
@(posedge clk);
#1;data_in = testData5[12052];
@(posedge clk);
#1;data_in = testData5[12053];
@(posedge clk);
#1;data_in = testData5[12054];
@(posedge clk);
#1;data_in = testData5[12055];
@(posedge clk);
#1;data_in = testData5[12056];
@(posedge clk);
#1;data_in = testData5[12057];
@(posedge clk);
#1;data_in = testData5[12058];
@(posedge clk);
#1;data_in = testData5[12059];
@(posedge clk);
#1;data_in = testData5[12060];
@(posedge clk);
#1;data_in = testData5[12061];
@(posedge clk);
#1;data_in = testData5[12062];
@(posedge clk);
#1;data_in = testData5[12063];
@(posedge clk);
#1;data_in = testData5[12064];
@(posedge clk);
#1;data_in = testData5[12065];
@(posedge clk);
#1;data_in = testData5[12066];
@(posedge clk);
#1;data_in = testData5[12067];
@(posedge clk);
#1;data_in = testData5[12068];
@(posedge clk);
#1;data_in = testData5[12069];
@(posedge clk);
#1;data_in = testData5[12070];
@(posedge clk);
#1;data_in = testData5[12071];
@(posedge clk);
#1;data_in = testData5[12072];
@(posedge clk);
#1;data_in = testData5[12073];
@(posedge clk);
#1;data_in = testData5[12074];
@(posedge clk);
#1;data_in = testData5[12075];
@(posedge clk);
#1;data_in = testData5[12076];
@(posedge clk);
#1;data_in = testData5[12077];
@(posedge clk);
#1;data_in = testData5[12078];
@(posedge clk);
#1;data_in = testData5[12079];
@(posedge clk);
#1;data_in = testData5[12080];
@(posedge clk);
#1;data_in = testData5[12081];
@(posedge clk);
#1;data_in = testData5[12082];
@(posedge clk);
#1;data_in = testData5[12083];
@(posedge clk);
#1;data_in = testData5[12084];
@(posedge clk);
#1;data_in = testData5[12085];
@(posedge clk);
#1;data_in = testData5[12086];
@(posedge clk);
#1;data_in = testData5[12087];
@(posedge clk);
#1;data_in = testData5[12088];
@(posedge clk);
#1;data_in = testData5[12089];
@(posedge clk);
#1;data_in = testData5[12090];
@(posedge clk);
#1;data_in = testData5[12091];
@(posedge clk);
#1;data_in = testData5[12092];
@(posedge clk);
#1;data_in = testData5[12093];
@(posedge clk);
#1;data_in = testData5[12094];
@(posedge clk);
#1;data_in = testData5[12095];
@(posedge clk);
#1;data_in = testData5[12096];
@(posedge clk);
#1;data_in = testData5[12097];
@(posedge clk);
#1;data_in = testData5[12098];
@(posedge clk);
#1;data_in = testData5[12099];
@(posedge clk);
#1;data_in = testData5[12100];
@(posedge clk);
#1;data_in = testData5[12101];
@(posedge clk);
#1;data_in = testData5[12102];
@(posedge clk);
#1;data_in = testData5[12103];
@(posedge clk);
#1;data_in = testData5[12104];
@(posedge clk);
#1;data_in = testData5[12105];
@(posedge clk);
#1;data_in = testData5[12106];
@(posedge clk);
#1;data_in = testData5[12107];
@(posedge clk);
#1;data_in = testData5[12108];
@(posedge clk);
#1;data_in = testData5[12109];
@(posedge clk);
#1;data_in = testData5[12110];
@(posedge clk);
#1;data_in = testData5[12111];
@(posedge clk);
#1;data_in = testData5[12112];
@(posedge clk);
#1;data_in = testData5[12113];
@(posedge clk);
#1;data_in = testData5[12114];
@(posedge clk);
#1;data_in = testData5[12115];
@(posedge clk);
#1;data_in = testData5[12116];
@(posedge clk);
#1;data_in = testData5[12117];
@(posedge clk);
#1;data_in = testData5[12118];
@(posedge clk);
#1;data_in = testData5[12119];
@(posedge clk);
#1;data_in = testData5[12120];
@(posedge clk);
#1;data_in = testData5[12121];
@(posedge clk);
#1;data_in = testData5[12122];
@(posedge clk);
#1;data_in = testData5[12123];
@(posedge clk);
#1;data_in = testData5[12124];
@(posedge clk);
#1;data_in = testData5[12125];
@(posedge clk);
#1;data_in = testData5[12126];
@(posedge clk);
#1;data_in = testData5[12127];
@(posedge clk);
#1;data_in = testData5[12128];
@(posedge clk);
#1;data_in = testData5[12129];
@(posedge clk);
#1;data_in = testData5[12130];
@(posedge clk);
#1;data_in = testData5[12131];
@(posedge clk);
#1;data_in = testData5[12132];
@(posedge clk);
#1;data_in = testData5[12133];
@(posedge clk);
#1;data_in = testData5[12134];
@(posedge clk);
#1;data_in = testData5[12135];
@(posedge clk);
#1;data_in = testData5[12136];
@(posedge clk);
#1;data_in = testData5[12137];
@(posedge clk);
#1;data_in = testData5[12138];
@(posedge clk);
#1;data_in = testData5[12139];
@(posedge clk);
#1;data_in = testData5[12140];
@(posedge clk);
#1;data_in = testData5[12141];
@(posedge clk);
#1;data_in = testData5[12142];
@(posedge clk);
#1;data_in = testData5[12143];
@(posedge clk);
#1;data_in = testData5[12144];
@(posedge clk);
#1;data_in = testData5[12145];
@(posedge clk);
#1;data_in = testData5[12146];
@(posedge clk);
#1;data_in = testData5[12147];
@(posedge clk);
#1;data_in = testData5[12148];
@(posedge clk);
#1;data_in = testData5[12149];
@(posedge clk);
#1;data_in = testData5[12150];
@(posedge clk);
#1;data_in = testData5[12151];
@(posedge clk);
#1;data_in = testData5[12152];
@(posedge clk);
#1;data_in = testData5[12153];
@(posedge clk);
#1;data_in = testData5[12154];
@(posedge clk);
#1;data_in = testData5[12155];
@(posedge clk);
#1;data_in = testData5[12156];
@(posedge clk);
#1;data_in = testData5[12157];
@(posedge clk);
#1;data_in = testData5[12158];
@(posedge clk);
#1;data_in = testData5[12159];
@(posedge clk);
#1;data_in = testData5[12160];
@(posedge clk);
#1;data_in = testData5[12161];
@(posedge clk);
#1;data_in = testData5[12162];
@(posedge clk);
#1;data_in = testData5[12163];
@(posedge clk);
#1;data_in = testData5[12164];
@(posedge clk);
#1;data_in = testData5[12165];
@(posedge clk);
#1;data_in = testData5[12166];
@(posedge clk);
#1;data_in = testData5[12167];
@(posedge clk);
#1;data_in = testData5[12168];
@(posedge clk);
#1;data_in = testData5[12169];
@(posedge clk);
#1;data_in = testData5[12170];
@(posedge clk);
#1;data_in = testData5[12171];
@(posedge clk);
#1;data_in = testData5[12172];
@(posedge clk);
#1;data_in = testData5[12173];
@(posedge clk);
#1;data_in = testData5[12174];
@(posedge clk);
#1;data_in = testData5[12175];
@(posedge clk);
#1;data_in = testData5[12176];
@(posedge clk);
#1;data_in = testData5[12177];
@(posedge clk);
#1;data_in = testData5[12178];
@(posedge clk);
#1;data_in = testData5[12179];
@(posedge clk);
#1;data_in = testData5[12180];
@(posedge clk);
#1;data_in = testData5[12181];
@(posedge clk);
#1;data_in = testData5[12182];
@(posedge clk);
#1;data_in = testData5[12183];
@(posedge clk);
#1;data_in = testData5[12184];
@(posedge clk);
#1;data_in = testData5[12185];
@(posedge clk);
#1;data_in = testData5[12186];
@(posedge clk);
#1;data_in = testData5[12187];
@(posedge clk);
#1;data_in = testData5[12188];
@(posedge clk);
#1;data_in = testData5[12189];
@(posedge clk);
#1;data_in = testData5[12190];
@(posedge clk);
#1;data_in = testData5[12191];
@(posedge clk);
#1;data_in = testData5[12192];
@(posedge clk);
#1;data_in = testData5[12193];
@(posedge clk);
#1;data_in = testData5[12194];
@(posedge clk);
#1;data_in = testData5[12195];
@(posedge clk);
#1;data_in = testData5[12196];
@(posedge clk);
#1;data_in = testData5[12197];
@(posedge clk);
#1;data_in = testData5[12198];
@(posedge clk);
#1;data_in = testData5[12199];
@(posedge clk);
#1;data_in = testData5[12200];
@(posedge clk);
#1;data_in = testData5[12201];
@(posedge clk);
#1;data_in = testData5[12202];
@(posedge clk);
#1;data_in = testData5[12203];
@(posedge clk);
#1;data_in = testData5[12204];
@(posedge clk);
#1;data_in = testData5[12205];
@(posedge clk);
#1;data_in = testData5[12206];
@(posedge clk);
#1;data_in = testData5[12207];
@(posedge clk);
#1;data_in = testData5[12208];
@(posedge clk);
#1;data_in = testData5[12209];
@(posedge clk);
#1;data_in = testData5[12210];
@(posedge clk);
#1;data_in = testData5[12211];
@(posedge clk);
#1;data_in = testData5[12212];
@(posedge clk);
#1;data_in = testData5[12213];
@(posedge clk);
#1;data_in = testData5[12214];
@(posedge clk);
#1;data_in = testData5[12215];
@(posedge clk);
#1;data_in = testData5[12216];
@(posedge clk);
#1;data_in = testData5[12217];
@(posedge clk);
#1;data_in = testData5[12218];
@(posedge clk);
#1;data_in = testData5[12219];
@(posedge clk);
#1;data_in = testData5[12220];
@(posedge clk);
#1;data_in = testData5[12221];
@(posedge clk);
#1;data_in = testData5[12222];
@(posedge clk);
#1;data_in = testData5[12223];
@(posedge clk);
#1;data_in = testData5[12224];
@(posedge clk);
#1;data_in = testData5[12225];
@(posedge clk);
#1;data_in = testData5[12226];
@(posedge clk);
#1;data_in = testData5[12227];
@(posedge clk);
#1;data_in = testData5[12228];
@(posedge clk);
#1;data_in = testData5[12229];
@(posedge clk);
#1;data_in = testData5[12230];
@(posedge clk);
#1;data_in = testData5[12231];
@(posedge clk);
#1;data_in = testData5[12232];
@(posedge clk);
#1;data_in = testData5[12233];
@(posedge clk);
#1;data_in = testData5[12234];
@(posedge clk);
#1;data_in = testData5[12235];
@(posedge clk);
#1;data_in = testData5[12236];
@(posedge clk);
#1;data_in = testData5[12237];
@(posedge clk);
#1;data_in = testData5[12238];
@(posedge clk);
#1;data_in = testData5[12239];
@(posedge clk);
#1;data_in = testData5[12240];
@(posedge clk);
#1;data_in = testData5[12241];
@(posedge clk);
#1;data_in = testData5[12242];
@(posedge clk);
#1;data_in = testData5[12243];
@(posedge clk);
#1;data_in = testData5[12244];
@(posedge clk);
#1;data_in = testData5[12245];
@(posedge clk);
#1;data_in = testData5[12246];
@(posedge clk);
#1;data_in = testData5[12247];
@(posedge clk);
#1;data_in = testData5[12248];
@(posedge clk);
#1;data_in = testData5[12249];
@(posedge clk);
#1;data_in = testData5[12250];
@(posedge clk);
#1;data_in = testData5[12251];
@(posedge clk);
#1;data_in = testData5[12252];
@(posedge clk);
#1;data_in = testData5[12253];
@(posedge clk);
#1;data_in = testData5[12254];
@(posedge clk);
#1;data_in = testData5[12255];
@(posedge clk);
#1;data_in = testData5[12256];
@(posedge clk);
#1;data_in = testData5[12257];
@(posedge clk);
#1;data_in = testData5[12258];
@(posedge clk);
#1;data_in = testData5[12259];
@(posedge clk);
#1;data_in = testData5[12260];
@(posedge clk);
#1;data_in = testData5[12261];
@(posedge clk);
#1;data_in = testData5[12262];
@(posedge clk);
#1;data_in = testData5[12263];
@(posedge clk);
#1;data_in = testData5[12264];
@(posedge clk);
#1;data_in = testData5[12265];
@(posedge clk);
#1;data_in = testData5[12266];
@(posedge clk);
#1;data_in = testData5[12267];
@(posedge clk);
#1;data_in = testData5[12268];
@(posedge clk);
#1;data_in = testData5[12269];
@(posedge clk);
#1;data_in = testData5[12270];
@(posedge clk);
#1;data_in = testData5[12271];
@(posedge clk);
#1;data_in = testData5[12272];
@(posedge clk);
#1;data_in = testData5[12273];
@(posedge clk);
#1;data_in = testData5[12274];
@(posedge clk);
#1;data_in = testData5[12275];
@(posedge clk);
#1;data_in = testData5[12276];
@(posedge clk);
#1;data_in = testData5[12277];
@(posedge clk);
#1;data_in = testData5[12278];
@(posedge clk);
#1;data_in = testData5[12279];
@(posedge clk);
#1;data_in = testData5[12280];
@(posedge clk);
#1;data_in = testData5[12281];
@(posedge clk);
#1;data_in = testData5[12282];
@(posedge clk);
#1;data_in = testData5[12283];
@(posedge clk);
#1;data_in = testData5[12284];
@(posedge clk);
#1;data_in = testData5[12285];
@(posedge clk);
#1;data_in = testData5[12286];
@(posedge clk);
#1;data_in = testData5[12287];
@(posedge clk);
#1;data_in = testData5[12288];
@(posedge clk);
#1;data_in = testData5[12289];
@(posedge clk);
#1;data_in = testData5[12290];
@(posedge clk);
#1;data_in = testData5[12291];
@(posedge clk);
#1;data_in = testData5[12292];
@(posedge clk);
#1;data_in = testData5[12293];
@(posedge clk);
#1;data_in = testData5[12294];
@(posedge clk);
#1;data_in = testData5[12295];
@(posedge clk);
#1;data_in = testData5[12296];
@(posedge clk);
#1;data_in = testData5[12297];
@(posedge clk);
#1;data_in = testData5[12298];
@(posedge clk);
#1;data_in = testData5[12299];
@(posedge clk);
#1;data_in = testData5[12300];
@(posedge clk);
#1;data_in = testData5[12301];
@(posedge clk);
#1;data_in = testData5[12302];
@(posedge clk);
#1;data_in = testData5[12303];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[12304]; 
@(posedge clk);
#1;data_in = testData5[12305];
@(posedge clk);
#1;data_in = testData5[12306];
@(posedge clk);
#1;data_in = testData5[12307];
@(posedge clk);
#1;data_in = testData5[12308];
@(posedge clk);
#1;data_in = testData5[12309];
@(posedge clk);
#1;data_in = testData5[12310];
@(posedge clk);
#1;data_in = testData5[12311];
@(posedge clk);
#1;data_in = testData5[12312];
@(posedge clk);
#1;data_in = testData5[12313];
@(posedge clk);
#1;data_in = testData5[12314];
@(posedge clk);
#1;data_in = testData5[12315];
@(posedge clk);
#1;data_in = testData5[12316];
@(posedge clk);
#1;data_in = testData5[12317];
@(posedge clk);
#1;data_in = testData5[12318];
@(posedge clk);
#1;data_in = testData5[12319];
@(posedge clk);
#1;data_in = testData5[12320];
@(posedge clk);
#1;data_in = testData5[12321];
@(posedge clk);
#1;data_in = testData5[12322];
@(posedge clk);
#1;data_in = testData5[12323];
@(posedge clk);
#1;data_in = testData5[12324];
@(posedge clk);
#1;data_in = testData5[12325];
@(posedge clk);
#1;data_in = testData5[12326];
@(posedge clk);
#1;data_in = testData5[12327];
@(posedge clk);
#1;data_in = testData5[12328];
@(posedge clk);
#1;data_in = testData5[12329];
@(posedge clk);
#1;data_in = testData5[12330];
@(posedge clk);
#1;data_in = testData5[12331];
@(posedge clk);
#1;data_in = testData5[12332];
@(posedge clk);
#1;data_in = testData5[12333];
@(posedge clk);
#1;data_in = testData5[12334];
@(posedge clk);
#1;data_in = testData5[12335];
@(posedge clk);
#1;data_in = testData5[12336];
@(posedge clk);
#1;data_in = testData5[12337];
@(posedge clk);
#1;data_in = testData5[12338];
@(posedge clk);
#1;data_in = testData5[12339];
@(posedge clk);
#1;data_in = testData5[12340];
@(posedge clk);
#1;data_in = testData5[12341];
@(posedge clk);
#1;data_in = testData5[12342];
@(posedge clk);
#1;data_in = testData5[12343];
@(posedge clk);
#1;data_in = testData5[12344];
@(posedge clk);
#1;data_in = testData5[12345];
@(posedge clk);
#1;data_in = testData5[12346];
@(posedge clk);
#1;data_in = testData5[12347];
@(posedge clk);
#1;data_in = testData5[12348];
@(posedge clk);
#1;data_in = testData5[12349];
@(posedge clk);
#1;data_in = testData5[12350];
@(posedge clk);
#1;data_in = testData5[12351];
@(posedge clk);
#1;data_in = testData5[12352];
@(posedge clk);
#1;data_in = testData5[12353];
@(posedge clk);
#1;data_in = testData5[12354];
@(posedge clk);
#1;data_in = testData5[12355];
@(posedge clk);
#1;data_in = testData5[12356];
@(posedge clk);
#1;data_in = testData5[12357];
@(posedge clk);
#1;data_in = testData5[12358];
@(posedge clk);
#1;data_in = testData5[12359];
@(posedge clk);
#1;data_in = testData5[12360];
@(posedge clk);
#1;data_in = testData5[12361];
@(posedge clk);
#1;data_in = testData5[12362];
@(posedge clk);
#1;data_in = testData5[12363];
@(posedge clk);
#1;data_in = testData5[12364];
@(posedge clk);
#1;data_in = testData5[12365];
@(posedge clk);
#1;data_in = testData5[12366];
@(posedge clk);
#1;data_in = testData5[12367];
@(posedge clk);
#1;data_in = testData5[12368];
@(posedge clk);
#1;data_in = testData5[12369];
@(posedge clk);
#1;data_in = testData5[12370];
@(posedge clk);
#1;data_in = testData5[12371];
@(posedge clk);
#1;data_in = testData5[12372];
@(posedge clk);
#1;data_in = testData5[12373];
@(posedge clk);
#1;data_in = testData5[12374];
@(posedge clk);
#1;data_in = testData5[12375];
@(posedge clk);
#1;data_in = testData5[12376];
@(posedge clk);
#1;data_in = testData5[12377];
@(posedge clk);
#1;data_in = testData5[12378];
@(posedge clk);
#1;data_in = testData5[12379];
@(posedge clk);
#1;data_in = testData5[12380];
@(posedge clk);
#1;data_in = testData5[12381];
@(posedge clk);
#1;data_in = testData5[12382];
@(posedge clk);
#1;data_in = testData5[12383];
@(posedge clk);
#1;data_in = testData5[12384];
@(posedge clk);
#1;data_in = testData5[12385];
@(posedge clk);
#1;data_in = testData5[12386];
@(posedge clk);
#1;data_in = testData5[12387];
@(posedge clk);
#1;data_in = testData5[12388];
@(posedge clk);
#1;data_in = testData5[12389];
@(posedge clk);
#1;data_in = testData5[12390];
@(posedge clk);
#1;data_in = testData5[12391];
@(posedge clk);
#1;data_in = testData5[12392];
@(posedge clk);
#1;data_in = testData5[12393];
@(posedge clk);
#1;data_in = testData5[12394];
@(posedge clk);
#1;data_in = testData5[12395];
@(posedge clk);
#1;data_in = testData5[12396];
@(posedge clk);
#1;data_in = testData5[12397];
@(posedge clk);
#1;data_in = testData5[12398];
@(posedge clk);
#1;data_in = testData5[12399];
@(posedge clk);
#1;data_in = testData5[12400];
@(posedge clk);
#1;data_in = testData5[12401];
@(posedge clk);
#1;data_in = testData5[12402];
@(posedge clk);
#1;data_in = testData5[12403];
@(posedge clk);
#1;data_in = testData5[12404];
@(posedge clk);
#1;data_in = testData5[12405];
@(posedge clk);
#1;data_in = testData5[12406];
@(posedge clk);
#1;data_in = testData5[12407];
@(posedge clk);
#1;data_in = testData5[12408];
@(posedge clk);
#1;data_in = testData5[12409];
@(posedge clk);
#1;data_in = testData5[12410];
@(posedge clk);
#1;data_in = testData5[12411];
@(posedge clk);
#1;data_in = testData5[12412];
@(posedge clk);
#1;data_in = testData5[12413];
@(posedge clk);
#1;data_in = testData5[12414];
@(posedge clk);
#1;data_in = testData5[12415];
@(posedge clk);
#1;data_in = testData5[12416];
@(posedge clk);
#1;data_in = testData5[12417];
@(posedge clk);
#1;data_in = testData5[12418];
@(posedge clk);
#1;data_in = testData5[12419];
@(posedge clk);
#1;data_in = testData5[12420];
@(posedge clk);
#1;data_in = testData5[12421];
@(posedge clk);
#1;data_in = testData5[12422];
@(posedge clk);
#1;data_in = testData5[12423];
@(posedge clk);
#1;data_in = testData5[12424];
@(posedge clk);
#1;data_in = testData5[12425];
@(posedge clk);
#1;data_in = testData5[12426];
@(posedge clk);
#1;data_in = testData5[12427];
@(posedge clk);
#1;data_in = testData5[12428];
@(posedge clk);
#1;data_in = testData5[12429];
@(posedge clk);
#1;data_in = testData5[12430];
@(posedge clk);
#1;data_in = testData5[12431];
@(posedge clk);
#1;data_in = testData5[12432];
@(posedge clk);
#1;data_in = testData5[12433];
@(posedge clk);
#1;data_in = testData5[12434];
@(posedge clk);
#1;data_in = testData5[12435];
@(posedge clk);
#1;data_in = testData5[12436];
@(posedge clk);
#1;data_in = testData5[12437];
@(posedge clk);
#1;data_in = testData5[12438];
@(posedge clk);
#1;data_in = testData5[12439];
@(posedge clk);
#1;data_in = testData5[12440];
@(posedge clk);
#1;data_in = testData5[12441];
@(posedge clk);
#1;data_in = testData5[12442];
@(posedge clk);
#1;data_in = testData5[12443];
@(posedge clk);
#1;data_in = testData5[12444];
@(posedge clk);
#1;data_in = testData5[12445];
@(posedge clk);
#1;data_in = testData5[12446];
@(posedge clk);
#1;data_in = testData5[12447];
@(posedge clk);
#1;data_in = testData5[12448];
@(posedge clk);
#1;data_in = testData5[12449];
@(posedge clk);
#1;data_in = testData5[12450];
@(posedge clk);
#1;data_in = testData5[12451];
@(posedge clk);
#1;data_in = testData5[12452];
@(posedge clk);
#1;data_in = testData5[12453];
@(posedge clk);
#1;data_in = testData5[12454];
@(posedge clk);
#1;data_in = testData5[12455];
@(posedge clk);
#1;data_in = testData5[12456];
@(posedge clk);
#1;data_in = testData5[12457];
@(posedge clk);
#1;data_in = testData5[12458];
@(posedge clk);
#1;data_in = testData5[12459];
@(posedge clk);
#1;data_in = testData5[12460];
@(posedge clk);
#1;data_in = testData5[12461];
@(posedge clk);
#1;data_in = testData5[12462];
@(posedge clk);
#1;data_in = testData5[12463];
@(posedge clk);
#1;data_in = testData5[12464];
@(posedge clk);
#1;data_in = testData5[12465];
@(posedge clk);
#1;data_in = testData5[12466];
@(posedge clk);
#1;data_in = testData5[12467];
@(posedge clk);
#1;data_in = testData5[12468];
@(posedge clk);
#1;data_in = testData5[12469];
@(posedge clk);
#1;data_in = testData5[12470];
@(posedge clk);
#1;data_in = testData5[12471];
@(posedge clk);
#1;data_in = testData5[12472];
@(posedge clk);
#1;data_in = testData5[12473];
@(posedge clk);
#1;data_in = testData5[12474];
@(posedge clk);
#1;data_in = testData5[12475];
@(posedge clk);
#1;data_in = testData5[12476];
@(posedge clk);
#1;data_in = testData5[12477];
@(posedge clk);
#1;data_in = testData5[12478];
@(posedge clk);
#1;data_in = testData5[12479];
@(posedge clk);
#1;data_in = testData5[12480];
@(posedge clk);
#1;data_in = testData5[12481];
@(posedge clk);
#1;data_in = testData5[12482];
@(posedge clk);
#1;data_in = testData5[12483];
@(posedge clk);
#1;data_in = testData5[12484];
@(posedge clk);
#1;data_in = testData5[12485];
@(posedge clk);
#1;data_in = testData5[12486];
@(posedge clk);
#1;data_in = testData5[12487];
@(posedge clk);
#1;data_in = testData5[12488];
@(posedge clk);
#1;data_in = testData5[12489];
@(posedge clk);
#1;data_in = testData5[12490];
@(posedge clk);
#1;data_in = testData5[12491];
@(posedge clk);
#1;data_in = testData5[12492];
@(posedge clk);
#1;data_in = testData5[12493];
@(posedge clk);
#1;data_in = testData5[12494];
@(posedge clk);
#1;data_in = testData5[12495];
@(posedge clk);
#1;data_in = testData5[12496];
@(posedge clk);
#1;data_in = testData5[12497];
@(posedge clk);
#1;data_in = testData5[12498];
@(posedge clk);
#1;data_in = testData5[12499];
@(posedge clk);
#1;data_in = testData5[12500];
@(posedge clk);
#1;data_in = testData5[12501];
@(posedge clk);
#1;data_in = testData5[12502];
@(posedge clk);
#1;data_in = testData5[12503];
@(posedge clk);
#1;data_in = testData5[12504];
@(posedge clk);
#1;data_in = testData5[12505];
@(posedge clk);
#1;data_in = testData5[12506];
@(posedge clk);
#1;data_in = testData5[12507];
@(posedge clk);
#1;data_in = testData5[12508];
@(posedge clk);
#1;data_in = testData5[12509];
@(posedge clk);
#1;data_in = testData5[12510];
@(posedge clk);
#1;data_in = testData5[12511];
@(posedge clk);
#1;data_in = testData5[12512];
@(posedge clk);
#1;data_in = testData5[12513];
@(posedge clk);
#1;data_in = testData5[12514];
@(posedge clk);
#1;data_in = testData5[12515];
@(posedge clk);
#1;data_in = testData5[12516];
@(posedge clk);
#1;data_in = testData5[12517];
@(posedge clk);
#1;data_in = testData5[12518];
@(posedge clk);
#1;data_in = testData5[12519];
@(posedge clk);
#1;data_in = testData5[12520];
@(posedge clk);
#1;data_in = testData5[12521];
@(posedge clk);
#1;data_in = testData5[12522];
@(posedge clk);
#1;data_in = testData5[12523];
@(posedge clk);
#1;data_in = testData5[12524];
@(posedge clk);
#1;data_in = testData5[12525];
@(posedge clk);
#1;data_in = testData5[12526];
@(posedge clk);
#1;data_in = testData5[12527];
@(posedge clk);
#1;data_in = testData5[12528];
@(posedge clk);
#1;data_in = testData5[12529];
@(posedge clk);
#1;data_in = testData5[12530];
@(posedge clk);
#1;data_in = testData5[12531];
@(posedge clk);
#1;data_in = testData5[12532];
@(posedge clk);
#1;data_in = testData5[12533];
@(posedge clk);
#1;data_in = testData5[12534];
@(posedge clk);
#1;data_in = testData5[12535];
@(posedge clk);
#1;data_in = testData5[12536];
@(posedge clk);
#1;data_in = testData5[12537];
@(posedge clk);
#1;data_in = testData5[12538];
@(posedge clk);
#1;data_in = testData5[12539];
@(posedge clk);
#1;data_in = testData5[12540];
@(posedge clk);
#1;data_in = testData5[12541];
@(posedge clk);
#1;data_in = testData5[12542];
@(posedge clk);
#1;data_in = testData5[12543];
@(posedge clk);
#1;data_in = testData5[12544];
@(posedge clk);
#1;data_in = testData5[12545];
@(posedge clk);
#1;data_in = testData5[12546];
@(posedge clk);
#1;data_in = testData5[12547];
@(posedge clk);
#1;data_in = testData5[12548];
@(posedge clk);
#1;data_in = testData5[12549];
@(posedge clk);
#1;data_in = testData5[12550];
@(posedge clk);
#1;data_in = testData5[12551];
@(posedge clk);
#1;data_in = testData5[12552];
@(posedge clk);
#1;data_in = testData5[12553];
@(posedge clk);
#1;data_in = testData5[12554];
@(posedge clk);
#1;data_in = testData5[12555];
@(posedge clk);
#1;data_in = testData5[12556];
@(posedge clk);
#1;data_in = testData5[12557];
@(posedge clk);
#1;data_in = testData5[12558];
@(posedge clk);
#1;data_in = testData5[12559];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[12560]; 
@(posedge clk);
#1;data_in = testData5[12561];
@(posedge clk);
#1;data_in = testData5[12562];
@(posedge clk);
#1;data_in = testData5[12563];
@(posedge clk);
#1;data_in = testData5[12564];
@(posedge clk);
#1;data_in = testData5[12565];
@(posedge clk);
#1;data_in = testData5[12566];
@(posedge clk);
#1;data_in = testData5[12567];
@(posedge clk);
#1;data_in = testData5[12568];
@(posedge clk);
#1;data_in = testData5[12569];
@(posedge clk);
#1;data_in = testData5[12570];
@(posedge clk);
#1;data_in = testData5[12571];
@(posedge clk);
#1;data_in = testData5[12572];
@(posedge clk);
#1;data_in = testData5[12573];
@(posedge clk);
#1;data_in = testData5[12574];
@(posedge clk);
#1;data_in = testData5[12575];
@(posedge clk);
#1;data_in = testData5[12576];
@(posedge clk);
#1;data_in = testData5[12577];
@(posedge clk);
#1;data_in = testData5[12578];
@(posedge clk);
#1;data_in = testData5[12579];
@(posedge clk);
#1;data_in = testData5[12580];
@(posedge clk);
#1;data_in = testData5[12581];
@(posedge clk);
#1;data_in = testData5[12582];
@(posedge clk);
#1;data_in = testData5[12583];
@(posedge clk);
#1;data_in = testData5[12584];
@(posedge clk);
#1;data_in = testData5[12585];
@(posedge clk);
#1;data_in = testData5[12586];
@(posedge clk);
#1;data_in = testData5[12587];
@(posedge clk);
#1;data_in = testData5[12588];
@(posedge clk);
#1;data_in = testData5[12589];
@(posedge clk);
#1;data_in = testData5[12590];
@(posedge clk);
#1;data_in = testData5[12591];
@(posedge clk);
#1;data_in = testData5[12592];
@(posedge clk);
#1;data_in = testData5[12593];
@(posedge clk);
#1;data_in = testData5[12594];
@(posedge clk);
#1;data_in = testData5[12595];
@(posedge clk);
#1;data_in = testData5[12596];
@(posedge clk);
#1;data_in = testData5[12597];
@(posedge clk);
#1;data_in = testData5[12598];
@(posedge clk);
#1;data_in = testData5[12599];
@(posedge clk);
#1;data_in = testData5[12600];
@(posedge clk);
#1;data_in = testData5[12601];
@(posedge clk);
#1;data_in = testData5[12602];
@(posedge clk);
#1;data_in = testData5[12603];
@(posedge clk);
#1;data_in = testData5[12604];
@(posedge clk);
#1;data_in = testData5[12605];
@(posedge clk);
#1;data_in = testData5[12606];
@(posedge clk);
#1;data_in = testData5[12607];
@(posedge clk);
#1;data_in = testData5[12608];
@(posedge clk);
#1;data_in = testData5[12609];
@(posedge clk);
#1;data_in = testData5[12610];
@(posedge clk);
#1;data_in = testData5[12611];
@(posedge clk);
#1;data_in = testData5[12612];
@(posedge clk);
#1;data_in = testData5[12613];
@(posedge clk);
#1;data_in = testData5[12614];
@(posedge clk);
#1;data_in = testData5[12615];
@(posedge clk);
#1;data_in = testData5[12616];
@(posedge clk);
#1;data_in = testData5[12617];
@(posedge clk);
#1;data_in = testData5[12618];
@(posedge clk);
#1;data_in = testData5[12619];
@(posedge clk);
#1;data_in = testData5[12620];
@(posedge clk);
#1;data_in = testData5[12621];
@(posedge clk);
#1;data_in = testData5[12622];
@(posedge clk);
#1;data_in = testData5[12623];
@(posedge clk);
#1;data_in = testData5[12624];
@(posedge clk);
#1;data_in = testData5[12625];
@(posedge clk);
#1;data_in = testData5[12626];
@(posedge clk);
#1;data_in = testData5[12627];
@(posedge clk);
#1;data_in = testData5[12628];
@(posedge clk);
#1;data_in = testData5[12629];
@(posedge clk);
#1;data_in = testData5[12630];
@(posedge clk);
#1;data_in = testData5[12631];
@(posedge clk);
#1;data_in = testData5[12632];
@(posedge clk);
#1;data_in = testData5[12633];
@(posedge clk);
#1;data_in = testData5[12634];
@(posedge clk);
#1;data_in = testData5[12635];
@(posedge clk);
#1;data_in = testData5[12636];
@(posedge clk);
#1;data_in = testData5[12637];
@(posedge clk);
#1;data_in = testData5[12638];
@(posedge clk);
#1;data_in = testData5[12639];
@(posedge clk);
#1;data_in = testData5[12640];
@(posedge clk);
#1;data_in = testData5[12641];
@(posedge clk);
#1;data_in = testData5[12642];
@(posedge clk);
#1;data_in = testData5[12643];
@(posedge clk);
#1;data_in = testData5[12644];
@(posedge clk);
#1;data_in = testData5[12645];
@(posedge clk);
#1;data_in = testData5[12646];
@(posedge clk);
#1;data_in = testData5[12647];
@(posedge clk);
#1;data_in = testData5[12648];
@(posedge clk);
#1;data_in = testData5[12649];
@(posedge clk);
#1;data_in = testData5[12650];
@(posedge clk);
#1;data_in = testData5[12651];
@(posedge clk);
#1;data_in = testData5[12652];
@(posedge clk);
#1;data_in = testData5[12653];
@(posedge clk);
#1;data_in = testData5[12654];
@(posedge clk);
#1;data_in = testData5[12655];
@(posedge clk);
#1;data_in = testData5[12656];
@(posedge clk);
#1;data_in = testData5[12657];
@(posedge clk);
#1;data_in = testData5[12658];
@(posedge clk);
#1;data_in = testData5[12659];
@(posedge clk);
#1;data_in = testData5[12660];
@(posedge clk);
#1;data_in = testData5[12661];
@(posedge clk);
#1;data_in = testData5[12662];
@(posedge clk);
#1;data_in = testData5[12663];
@(posedge clk);
#1;data_in = testData5[12664];
@(posedge clk);
#1;data_in = testData5[12665];
@(posedge clk);
#1;data_in = testData5[12666];
@(posedge clk);
#1;data_in = testData5[12667];
@(posedge clk);
#1;data_in = testData5[12668];
@(posedge clk);
#1;data_in = testData5[12669];
@(posedge clk);
#1;data_in = testData5[12670];
@(posedge clk);
#1;data_in = testData5[12671];
@(posedge clk);
#1;data_in = testData5[12672];
@(posedge clk);
#1;data_in = testData5[12673];
@(posedge clk);
#1;data_in = testData5[12674];
@(posedge clk);
#1;data_in = testData5[12675];
@(posedge clk);
#1;data_in = testData5[12676];
@(posedge clk);
#1;data_in = testData5[12677];
@(posedge clk);
#1;data_in = testData5[12678];
@(posedge clk);
#1;data_in = testData5[12679];
@(posedge clk);
#1;data_in = testData5[12680];
@(posedge clk);
#1;data_in = testData5[12681];
@(posedge clk);
#1;data_in = testData5[12682];
@(posedge clk);
#1;data_in = testData5[12683];
@(posedge clk);
#1;data_in = testData5[12684];
@(posedge clk);
#1;data_in = testData5[12685];
@(posedge clk);
#1;data_in = testData5[12686];
@(posedge clk);
#1;data_in = testData5[12687];
@(posedge clk);
#1;data_in = testData5[12688];
@(posedge clk);
#1;data_in = testData5[12689];
@(posedge clk);
#1;data_in = testData5[12690];
@(posedge clk);
#1;data_in = testData5[12691];
@(posedge clk);
#1;data_in = testData5[12692];
@(posedge clk);
#1;data_in = testData5[12693];
@(posedge clk);
#1;data_in = testData5[12694];
@(posedge clk);
#1;data_in = testData5[12695];
@(posedge clk);
#1;data_in = testData5[12696];
@(posedge clk);
#1;data_in = testData5[12697];
@(posedge clk);
#1;data_in = testData5[12698];
@(posedge clk);
#1;data_in = testData5[12699];
@(posedge clk);
#1;data_in = testData5[12700];
@(posedge clk);
#1;data_in = testData5[12701];
@(posedge clk);
#1;data_in = testData5[12702];
@(posedge clk);
#1;data_in = testData5[12703];
@(posedge clk);
#1;data_in = testData5[12704];
@(posedge clk);
#1;data_in = testData5[12705];
@(posedge clk);
#1;data_in = testData5[12706];
@(posedge clk);
#1;data_in = testData5[12707];
@(posedge clk);
#1;data_in = testData5[12708];
@(posedge clk);
#1;data_in = testData5[12709];
@(posedge clk);
#1;data_in = testData5[12710];
@(posedge clk);
#1;data_in = testData5[12711];
@(posedge clk);
#1;data_in = testData5[12712];
@(posedge clk);
#1;data_in = testData5[12713];
@(posedge clk);
#1;data_in = testData5[12714];
@(posedge clk);
#1;data_in = testData5[12715];
@(posedge clk);
#1;data_in = testData5[12716];
@(posedge clk);
#1;data_in = testData5[12717];
@(posedge clk);
#1;data_in = testData5[12718];
@(posedge clk);
#1;data_in = testData5[12719];
@(posedge clk);
#1;data_in = testData5[12720];
@(posedge clk);
#1;data_in = testData5[12721];
@(posedge clk);
#1;data_in = testData5[12722];
@(posedge clk);
#1;data_in = testData5[12723];
@(posedge clk);
#1;data_in = testData5[12724];
@(posedge clk);
#1;data_in = testData5[12725];
@(posedge clk);
#1;data_in = testData5[12726];
@(posedge clk);
#1;data_in = testData5[12727];
@(posedge clk);
#1;data_in = testData5[12728];
@(posedge clk);
#1;data_in = testData5[12729];
@(posedge clk);
#1;data_in = testData5[12730];
@(posedge clk);
#1;data_in = testData5[12731];
@(posedge clk);
#1;data_in = testData5[12732];
@(posedge clk);
#1;data_in = testData5[12733];
@(posedge clk);
#1;data_in = testData5[12734];
@(posedge clk);
#1;data_in = testData5[12735];
@(posedge clk);
#1;data_in = testData5[12736];
@(posedge clk);
#1;data_in = testData5[12737];
@(posedge clk);
#1;data_in = testData5[12738];
@(posedge clk);
#1;data_in = testData5[12739];
@(posedge clk);
#1;data_in = testData5[12740];
@(posedge clk);
#1;data_in = testData5[12741];
@(posedge clk);
#1;data_in = testData5[12742];
@(posedge clk);
#1;data_in = testData5[12743];
@(posedge clk);
#1;data_in = testData5[12744];
@(posedge clk);
#1;data_in = testData5[12745];
@(posedge clk);
#1;data_in = testData5[12746];
@(posedge clk);
#1;data_in = testData5[12747];
@(posedge clk);
#1;data_in = testData5[12748];
@(posedge clk);
#1;data_in = testData5[12749];
@(posedge clk);
#1;data_in = testData5[12750];
@(posedge clk);
#1;data_in = testData5[12751];
@(posedge clk);
#1;data_in = testData5[12752];
@(posedge clk);
#1;data_in = testData5[12753];
@(posedge clk);
#1;data_in = testData5[12754];
@(posedge clk);
#1;data_in = testData5[12755];
@(posedge clk);
#1;data_in = testData5[12756];
@(posedge clk);
#1;data_in = testData5[12757];
@(posedge clk);
#1;data_in = testData5[12758];
@(posedge clk);
#1;data_in = testData5[12759];
@(posedge clk);
#1;data_in = testData5[12760];
@(posedge clk);
#1;data_in = testData5[12761];
@(posedge clk);
#1;data_in = testData5[12762];
@(posedge clk);
#1;data_in = testData5[12763];
@(posedge clk);
#1;data_in = testData5[12764];
@(posedge clk);
#1;data_in = testData5[12765];
@(posedge clk);
#1;data_in = testData5[12766];
@(posedge clk);
#1;data_in = testData5[12767];
@(posedge clk);
#1;data_in = testData5[12768];
@(posedge clk);
#1;data_in = testData5[12769];
@(posedge clk);
#1;data_in = testData5[12770];
@(posedge clk);
#1;data_in = testData5[12771];
@(posedge clk);
#1;data_in = testData5[12772];
@(posedge clk);
#1;data_in = testData5[12773];
@(posedge clk);
#1;data_in = testData5[12774];
@(posedge clk);
#1;data_in = testData5[12775];
@(posedge clk);
#1;data_in = testData5[12776];
@(posedge clk);
#1;data_in = testData5[12777];
@(posedge clk);
#1;data_in = testData5[12778];
@(posedge clk);
#1;data_in = testData5[12779];
@(posedge clk);
#1;data_in = testData5[12780];
@(posedge clk);
#1;data_in = testData5[12781];
@(posedge clk);
#1;data_in = testData5[12782];
@(posedge clk);
#1;data_in = testData5[12783];
@(posedge clk);
#1;data_in = testData5[12784];
@(posedge clk);
#1;data_in = testData5[12785];
@(posedge clk);
#1;data_in = testData5[12786];
@(posedge clk);
#1;data_in = testData5[12787];
@(posedge clk);
#1;data_in = testData5[12788];
@(posedge clk);
#1;data_in = testData5[12789];
@(posedge clk);
#1;data_in = testData5[12790];
@(posedge clk);
#1;data_in = testData5[12791];
@(posedge clk);
#1;data_in = testData5[12792];
@(posedge clk);
#1;data_in = testData5[12793];
@(posedge clk);
#1;data_in = testData5[12794];
@(posedge clk);
#1;data_in = testData5[12795];
@(posedge clk);
#1;data_in = testData5[12796];
@(posedge clk);
#1;data_in = testData5[12797];
@(posedge clk);
#1;data_in = testData5[12798];
@(posedge clk);
#1;data_in = testData5[12799];
@(posedge clk);
#1;data_in = testData5[12800];
@(posedge clk);
#1;data_in = testData5[12801];
@(posedge clk);
#1;data_in = testData5[12802];
@(posedge clk);
#1;data_in = testData5[12803];
@(posedge clk);
#1;data_in = testData5[12804];
@(posedge clk);
#1;data_in = testData5[12805];
@(posedge clk);
#1;data_in = testData5[12806];
@(posedge clk);
#1;data_in = testData5[12807];
@(posedge clk);
#1;data_in = testData5[12808];
@(posedge clk);
#1;data_in = testData5[12809];
@(posedge clk);
#1;data_in = testData5[12810];
@(posedge clk);
#1;data_in = testData5[12811];
@(posedge clk);
#1;data_in = testData5[12812];
@(posedge clk);
#1;data_in = testData5[12813];
@(posedge clk);
#1;data_in = testData5[12814];
@(posedge clk);
#1;data_in = testData5[12815];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[12816]; 
@(posedge clk);
#1;data_in = testData5[12817];
@(posedge clk);
#1;data_in = testData5[12818];
@(posedge clk);
#1;data_in = testData5[12819];
@(posedge clk);
#1;data_in = testData5[12820];
@(posedge clk);
#1;data_in = testData5[12821];
@(posedge clk);
#1;data_in = testData5[12822];
@(posedge clk);
#1;data_in = testData5[12823];
@(posedge clk);
#1;data_in = testData5[12824];
@(posedge clk);
#1;data_in = testData5[12825];
@(posedge clk);
#1;data_in = testData5[12826];
@(posedge clk);
#1;data_in = testData5[12827];
@(posedge clk);
#1;data_in = testData5[12828];
@(posedge clk);
#1;data_in = testData5[12829];
@(posedge clk);
#1;data_in = testData5[12830];
@(posedge clk);
#1;data_in = testData5[12831];
@(posedge clk);
#1;data_in = testData5[12832];
@(posedge clk);
#1;data_in = testData5[12833];
@(posedge clk);
#1;data_in = testData5[12834];
@(posedge clk);
#1;data_in = testData5[12835];
@(posedge clk);
#1;data_in = testData5[12836];
@(posedge clk);
#1;data_in = testData5[12837];
@(posedge clk);
#1;data_in = testData5[12838];
@(posedge clk);
#1;data_in = testData5[12839];
@(posedge clk);
#1;data_in = testData5[12840];
@(posedge clk);
#1;data_in = testData5[12841];
@(posedge clk);
#1;data_in = testData5[12842];
@(posedge clk);
#1;data_in = testData5[12843];
@(posedge clk);
#1;data_in = testData5[12844];
@(posedge clk);
#1;data_in = testData5[12845];
@(posedge clk);
#1;data_in = testData5[12846];
@(posedge clk);
#1;data_in = testData5[12847];
@(posedge clk);
#1;data_in = testData5[12848];
@(posedge clk);
#1;data_in = testData5[12849];
@(posedge clk);
#1;data_in = testData5[12850];
@(posedge clk);
#1;data_in = testData5[12851];
@(posedge clk);
#1;data_in = testData5[12852];
@(posedge clk);
#1;data_in = testData5[12853];
@(posedge clk);
#1;data_in = testData5[12854];
@(posedge clk);
#1;data_in = testData5[12855];
@(posedge clk);
#1;data_in = testData5[12856];
@(posedge clk);
#1;data_in = testData5[12857];
@(posedge clk);
#1;data_in = testData5[12858];
@(posedge clk);
#1;data_in = testData5[12859];
@(posedge clk);
#1;data_in = testData5[12860];
@(posedge clk);
#1;data_in = testData5[12861];
@(posedge clk);
#1;data_in = testData5[12862];
@(posedge clk);
#1;data_in = testData5[12863];
@(posedge clk);
#1;data_in = testData5[12864];
@(posedge clk);
#1;data_in = testData5[12865];
@(posedge clk);
#1;data_in = testData5[12866];
@(posedge clk);
#1;data_in = testData5[12867];
@(posedge clk);
#1;data_in = testData5[12868];
@(posedge clk);
#1;data_in = testData5[12869];
@(posedge clk);
#1;data_in = testData5[12870];
@(posedge clk);
#1;data_in = testData5[12871];
@(posedge clk);
#1;data_in = testData5[12872];
@(posedge clk);
#1;data_in = testData5[12873];
@(posedge clk);
#1;data_in = testData5[12874];
@(posedge clk);
#1;data_in = testData5[12875];
@(posedge clk);
#1;data_in = testData5[12876];
@(posedge clk);
#1;data_in = testData5[12877];
@(posedge clk);
#1;data_in = testData5[12878];
@(posedge clk);
#1;data_in = testData5[12879];
@(posedge clk);
#1;data_in = testData5[12880];
@(posedge clk);
#1;data_in = testData5[12881];
@(posedge clk);
#1;data_in = testData5[12882];
@(posedge clk);
#1;data_in = testData5[12883];
@(posedge clk);
#1;data_in = testData5[12884];
@(posedge clk);
#1;data_in = testData5[12885];
@(posedge clk);
#1;data_in = testData5[12886];
@(posedge clk);
#1;data_in = testData5[12887];
@(posedge clk);
#1;data_in = testData5[12888];
@(posedge clk);
#1;data_in = testData5[12889];
@(posedge clk);
#1;data_in = testData5[12890];
@(posedge clk);
#1;data_in = testData5[12891];
@(posedge clk);
#1;data_in = testData5[12892];
@(posedge clk);
#1;data_in = testData5[12893];
@(posedge clk);
#1;data_in = testData5[12894];
@(posedge clk);
#1;data_in = testData5[12895];
@(posedge clk);
#1;data_in = testData5[12896];
@(posedge clk);
#1;data_in = testData5[12897];
@(posedge clk);
#1;data_in = testData5[12898];
@(posedge clk);
#1;data_in = testData5[12899];
@(posedge clk);
#1;data_in = testData5[12900];
@(posedge clk);
#1;data_in = testData5[12901];
@(posedge clk);
#1;data_in = testData5[12902];
@(posedge clk);
#1;data_in = testData5[12903];
@(posedge clk);
#1;data_in = testData5[12904];
@(posedge clk);
#1;data_in = testData5[12905];
@(posedge clk);
#1;data_in = testData5[12906];
@(posedge clk);
#1;data_in = testData5[12907];
@(posedge clk);
#1;data_in = testData5[12908];
@(posedge clk);
#1;data_in = testData5[12909];
@(posedge clk);
#1;data_in = testData5[12910];
@(posedge clk);
#1;data_in = testData5[12911];
@(posedge clk);
#1;data_in = testData5[12912];
@(posedge clk);
#1;data_in = testData5[12913];
@(posedge clk);
#1;data_in = testData5[12914];
@(posedge clk);
#1;data_in = testData5[12915];
@(posedge clk);
#1;data_in = testData5[12916];
@(posedge clk);
#1;data_in = testData5[12917];
@(posedge clk);
#1;data_in = testData5[12918];
@(posedge clk);
#1;data_in = testData5[12919];
@(posedge clk);
#1;data_in = testData5[12920];
@(posedge clk);
#1;data_in = testData5[12921];
@(posedge clk);
#1;data_in = testData5[12922];
@(posedge clk);
#1;data_in = testData5[12923];
@(posedge clk);
#1;data_in = testData5[12924];
@(posedge clk);
#1;data_in = testData5[12925];
@(posedge clk);
#1;data_in = testData5[12926];
@(posedge clk);
#1;data_in = testData5[12927];
@(posedge clk);
#1;data_in = testData5[12928];
@(posedge clk);
#1;data_in = testData5[12929];
@(posedge clk);
#1;data_in = testData5[12930];
@(posedge clk);
#1;data_in = testData5[12931];
@(posedge clk);
#1;data_in = testData5[12932];
@(posedge clk);
#1;data_in = testData5[12933];
@(posedge clk);
#1;data_in = testData5[12934];
@(posedge clk);
#1;data_in = testData5[12935];
@(posedge clk);
#1;data_in = testData5[12936];
@(posedge clk);
#1;data_in = testData5[12937];
@(posedge clk);
#1;data_in = testData5[12938];
@(posedge clk);
#1;data_in = testData5[12939];
@(posedge clk);
#1;data_in = testData5[12940];
@(posedge clk);
#1;data_in = testData5[12941];
@(posedge clk);
#1;data_in = testData5[12942];
@(posedge clk);
#1;data_in = testData5[12943];
@(posedge clk);
#1;data_in = testData5[12944];
@(posedge clk);
#1;data_in = testData5[12945];
@(posedge clk);
#1;data_in = testData5[12946];
@(posedge clk);
#1;data_in = testData5[12947];
@(posedge clk);
#1;data_in = testData5[12948];
@(posedge clk);
#1;data_in = testData5[12949];
@(posedge clk);
#1;data_in = testData5[12950];
@(posedge clk);
#1;data_in = testData5[12951];
@(posedge clk);
#1;data_in = testData5[12952];
@(posedge clk);
#1;data_in = testData5[12953];
@(posedge clk);
#1;data_in = testData5[12954];
@(posedge clk);
#1;data_in = testData5[12955];
@(posedge clk);
#1;data_in = testData5[12956];
@(posedge clk);
#1;data_in = testData5[12957];
@(posedge clk);
#1;data_in = testData5[12958];
@(posedge clk);
#1;data_in = testData5[12959];
@(posedge clk);
#1;data_in = testData5[12960];
@(posedge clk);
#1;data_in = testData5[12961];
@(posedge clk);
#1;data_in = testData5[12962];
@(posedge clk);
#1;data_in = testData5[12963];
@(posedge clk);
#1;data_in = testData5[12964];
@(posedge clk);
#1;data_in = testData5[12965];
@(posedge clk);
#1;data_in = testData5[12966];
@(posedge clk);
#1;data_in = testData5[12967];
@(posedge clk);
#1;data_in = testData5[12968];
@(posedge clk);
#1;data_in = testData5[12969];
@(posedge clk);
#1;data_in = testData5[12970];
@(posedge clk);
#1;data_in = testData5[12971];
@(posedge clk);
#1;data_in = testData5[12972];
@(posedge clk);
#1;data_in = testData5[12973];
@(posedge clk);
#1;data_in = testData5[12974];
@(posedge clk);
#1;data_in = testData5[12975];
@(posedge clk);
#1;data_in = testData5[12976];
@(posedge clk);
#1;data_in = testData5[12977];
@(posedge clk);
#1;data_in = testData5[12978];
@(posedge clk);
#1;data_in = testData5[12979];
@(posedge clk);
#1;data_in = testData5[12980];
@(posedge clk);
#1;data_in = testData5[12981];
@(posedge clk);
#1;data_in = testData5[12982];
@(posedge clk);
#1;data_in = testData5[12983];
@(posedge clk);
#1;data_in = testData5[12984];
@(posedge clk);
#1;data_in = testData5[12985];
@(posedge clk);
#1;data_in = testData5[12986];
@(posedge clk);
#1;data_in = testData5[12987];
@(posedge clk);
#1;data_in = testData5[12988];
@(posedge clk);
#1;data_in = testData5[12989];
@(posedge clk);
#1;data_in = testData5[12990];
@(posedge clk);
#1;data_in = testData5[12991];
@(posedge clk);
#1;data_in = testData5[12992];
@(posedge clk);
#1;data_in = testData5[12993];
@(posedge clk);
#1;data_in = testData5[12994];
@(posedge clk);
#1;data_in = testData5[12995];
@(posedge clk);
#1;data_in = testData5[12996];
@(posedge clk);
#1;data_in = testData5[12997];
@(posedge clk);
#1;data_in = testData5[12998];
@(posedge clk);
#1;data_in = testData5[12999];
@(posedge clk);
#1;data_in = testData5[13000];
@(posedge clk);
#1;data_in = testData5[13001];
@(posedge clk);
#1;data_in = testData5[13002];
@(posedge clk);
#1;data_in = testData5[13003];
@(posedge clk);
#1;data_in = testData5[13004];
@(posedge clk);
#1;data_in = testData5[13005];
@(posedge clk);
#1;data_in = testData5[13006];
@(posedge clk);
#1;data_in = testData5[13007];
@(posedge clk);
#1;data_in = testData5[13008];
@(posedge clk);
#1;data_in = testData5[13009];
@(posedge clk);
#1;data_in = testData5[13010];
@(posedge clk);
#1;data_in = testData5[13011];
@(posedge clk);
#1;data_in = testData5[13012];
@(posedge clk);
#1;data_in = testData5[13013];
@(posedge clk);
#1;data_in = testData5[13014];
@(posedge clk);
#1;data_in = testData5[13015];
@(posedge clk);
#1;data_in = testData5[13016];
@(posedge clk);
#1;data_in = testData5[13017];
@(posedge clk);
#1;data_in = testData5[13018];
@(posedge clk);
#1;data_in = testData5[13019];
@(posedge clk);
#1;data_in = testData5[13020];
@(posedge clk);
#1;data_in = testData5[13021];
@(posedge clk);
#1;data_in = testData5[13022];
@(posedge clk);
#1;data_in = testData5[13023];
@(posedge clk);
#1;data_in = testData5[13024];
@(posedge clk);
#1;data_in = testData5[13025];
@(posedge clk);
#1;data_in = testData5[13026];
@(posedge clk);
#1;data_in = testData5[13027];
@(posedge clk);
#1;data_in = testData5[13028];
@(posedge clk);
#1;data_in = testData5[13029];
@(posedge clk);
#1;data_in = testData5[13030];
@(posedge clk);
#1;data_in = testData5[13031];
@(posedge clk);
#1;data_in = testData5[13032];
@(posedge clk);
#1;data_in = testData5[13033];
@(posedge clk);
#1;data_in = testData5[13034];
@(posedge clk);
#1;data_in = testData5[13035];
@(posedge clk);
#1;data_in = testData5[13036];
@(posedge clk);
#1;data_in = testData5[13037];
@(posedge clk);
#1;data_in = testData5[13038];
@(posedge clk);
#1;data_in = testData5[13039];
@(posedge clk);
#1;data_in = testData5[13040];
@(posedge clk);
#1;data_in = testData5[13041];
@(posedge clk);
#1;data_in = testData5[13042];
@(posedge clk);
#1;data_in = testData5[13043];
@(posedge clk);
#1;data_in = testData5[13044];
@(posedge clk);
#1;data_in = testData5[13045];
@(posedge clk);
#1;data_in = testData5[13046];
@(posedge clk);
#1;data_in = testData5[13047];
@(posedge clk);
#1;data_in = testData5[13048];
@(posedge clk);
#1;data_in = testData5[13049];
@(posedge clk);
#1;data_in = testData5[13050];
@(posedge clk);
#1;data_in = testData5[13051];
@(posedge clk);
#1;data_in = testData5[13052];
@(posedge clk);
#1;data_in = testData5[13053];
@(posedge clk);
#1;data_in = testData5[13054];
@(posedge clk);
#1;data_in = testData5[13055];
@(posedge clk);
#1;data_in = testData5[13056];
@(posedge clk);
#1;data_in = testData5[13057];
@(posedge clk);
#1;data_in = testData5[13058];
@(posedge clk);
#1;data_in = testData5[13059];
@(posedge clk);
#1;data_in = testData5[13060];
@(posedge clk);
#1;data_in = testData5[13061];
@(posedge clk);
#1;data_in = testData5[13062];
@(posedge clk);
#1;data_in = testData5[13063];
@(posedge clk);
#1;data_in = testData5[13064];
@(posedge clk);
#1;data_in = testData5[13065];
@(posedge clk);
#1;data_in = testData5[13066];
@(posedge clk);
#1;data_in = testData5[13067];
@(posedge clk);
#1;data_in = testData5[13068];
@(posedge clk);
#1;data_in = testData5[13069];
@(posedge clk);
#1;data_in = testData5[13070];
@(posedge clk);
#1;data_in = testData5[13071];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[8] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[9] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[10] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[11] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[12] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[13] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[14] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[15] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
